`ifndef DEFINES_H_
`define DEFINES_H_

`define ALU_OPW 7

`define ALU_OP_ADD 0
`define ALU_OP_SUB 1
`define ALU_OP_AND 2
`define ALU_OP_OR 3
`define ALU_OP_XOR 4
`define ALU_OP_SLL 5
`define ALU_OP_SRL 6

`endif
