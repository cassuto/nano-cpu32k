// GaoZiBo

module mycpu(
   input clk,
   input rst_n
);

   

endmodule