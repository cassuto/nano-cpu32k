/*
Copyright 2021 GaoZiBo <diyer175@hotmail.com>
Powered by YSYX https://oscpu.github.io/ysyx

Licensed under The MIT License (MIT).
-------------------------------------
Permission is hereby granted, free of charge, to any person obtaining a copy of
this software and associated documentation files (the "Software"), to deal in
the Software without restriction, including without limitation the rights to
use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of
the Software, and to permit persons to whom the Software is furnished to do so,
subject to the following conditions:

The above copyright notice and this permission notice shall be included in all
copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED,INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, FITNESS
FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR
COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER
IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 */

`include "ncpu64k_config.vh"

module ifu
#(
   parameter CONFIG_AW = 0,
   parameter CONFIG_P_FETCH_WIDTH = 0,
   parameter CONFIG_P_ISSUE_WIDTH = 0,
   parameter CONFIG_P_IQ_DEPTH = 0,
   parameter CONFIG_P_PAGE_SIZE = 0,
   parameter CONFIG_IC_P_LINE = 0,
   parameter CONFIG_IC_P_SETS = 0,
   parameter CONFIG_IC_P_WAYS = 0,
   parameter CONFIG_PHT_P_NUM = 0,
   parameter CONFIG_BTB_P_NUM = 0,
   parameter AXI_P_DW_BYTES = 0,
   parameter AXI_ADDR_WIDTH = 0,
   parameter AXI_ID_WIDTH = 0,
   parameter AXI_USER_WIDTH = 0
)
(
   input                               clk,
   input                               rst,
   input                               flush,
   input [CONFIG_AW-1:0]               flush_tgt,
   // To ID
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_valid,
   input [CONFIG_P_ISSUE_WIDTH:0]      id_pop_cnt,
   output [`NCPU_INSN_DW * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_ins,
   output [CONFIG_AW * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_pc,
   output [`FNT_EXC_W * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_exc,
   output [`BPU_UPD_W*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_bpu_upd,
   // From EX
   input                               icop_inv,
   input [CONFIG_AW-1:0]               icop_inv_paddr,
   input                               bpu_wb,
   input                               bpu_wb_is_bcc,
   input                               bpu_wb_is_breg,
   input                               bpu_wb_bcc_taken,
   input [CONFIG_AW-3:0]               bpu_wb_pc,
   input [CONFIG_AW-3:0]               bpu_wb_npc_act,
   input [`BPU_UPD_W-1:0]              bpu_wb_upd,
   // To EX
   output                              icop_stall_req,
   // AXI Master
   input                               axi_ar_ready_i,
   output                              axi_ar_valid_o,
   output [AXI_ADDR_WIDTH-1:0]         axi_ar_addr_o,
   output [2:0]                        axi_ar_prot_o,
   output [AXI_ID_WIDTH-1:0]           axi_ar_id_o,
   output [AXI_USER_WIDTH-1:0]         axi_ar_user_o,
   output [7:0]                        axi_ar_len_o,
   output [2:0]                        axi_ar_size_o,
   output [1:0]                        axi_ar_burst_o,
   output                              axi_ar_lock_o,
   output [3:0]                        axi_ar_cache_o,
   output [3:0]                        axi_ar_qos_o,
   output [3:0]                        axi_ar_region_o,

   output                              axi_r_ready_o,
   input                               axi_r_valid_i,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  axi_r_data_i,
   input  [1:0]                        axi_r_resp_i,
   input                               axi_r_last_i,
   input  [AXI_ID_WIDTH-1:0]           axi_r_id_i,
   input  [AXI_USER_WIDTH-1:0]         axi_r_user_i
);
   localparam P_FETCH_DW_BYTES         = (`NCPU_P_INSN_LEN + CONFIG_P_FETCH_WIDTH);
   localparam FW                       = (1<<CONFIG_P_FETCH_WIDTH);
   
   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire                 ic_stall_req;           // From U_ICACHE of icache.v
   wire                 iq_ready;               // From U_IQ of iq.v
   // End of automatics
   wire                                p_ce;
   wire [CONFIG_P_PAGE_SIZE-1:0]       vpo;
   wire [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] ppn_s2;
   wire                                kill_req_s2;
   wire                                pred_branch_taken;
   wire [CONFIG_AW-1:0]                pc;
   reg [CONFIG_AW-1:0]                 pc_nxt;
   // Stage 1 Input
   wire [CONFIG_AW-1:0]                s1i_fetch_vaddr;
   wire [FW-1:0]                       s1i_fetch_valid;
   reg [FW-1:0]                        s1i_valid_msk;
   wire [CONFIG_AW-1:0]                s1i_pc                           [FW-1:0];
   wire [(CONFIG_AW-2)*FW-1:0]         s1i_bpu_pc;
   wire [CONFIG_P_FETCH_WIDTH:0]       s1i_push_cnt;
   // Stage 2 Input / Stage 1 Output
   wire [CONFIG_AW-1:0]                s1o_pc                           [FW-1:0];
   wire [`FNT_EXC_W-1:0]               s1o_exc;
   wire [CONFIG_P_FETCH_WIDTH:0]       s1o_push_cnt;
   wire [(CONFIG_AW-2)*FW-1:0]         s1o_bpu_npc_packed;
   wire [CONFIG_AW-3:0]                s1o_bpu_npc                      [FW-1:0];
   wire [`BPU_UPD_W*FW-1:0]            s1o_bpu_upd_packed;
   wire [`BPU_UPD_W-1:0]               s1o_bpu_upd                      [FW-1:0];
   wire [FW-1:0]                       s1o_bpu_taken;
   wire [CONFIG_P_FETCH_WIDTH-1:0]     s1o_bpu_taken_inst_idx;
   wire [`BPU_UPD_W-1:0]               s2i_bpu_upd                      [FW-1:0];
   // Stage 3 Input / Stage 2 Output
   wire [CONFIG_AW-1:0]                s2o_pc                           [FW-1:0];
   wire [`FNT_EXC_W-1:0]               s2o_exc;
   wire [`BPU_UPD_W-1:0]               s2o_bpu_upd                      [FW-1:0];
   wire                                s2o_valid;
   wire [CONFIG_P_FETCH_WIDTH:0]       s2o_push_cnt;
   wire [`NCPU_INSN_DW*FW-1:0]         iq_ins;
   wire [CONFIG_AW*FW-1:0]             iq_pc;
   wire [`FNT_EXC_W*FW-1:0]            iq_exc;
   wire [`BPU_UPD_W*FW-1:0]            iq_bpu_upd;
   wire [CONFIG_P_FETCH_WIDTH:0]       iq_push_cnt;
   
   genvar i;
   integer j;

/* icache AUTO_TEMPLATE (
      .stall_req                       (ic_stall_req),
      .ins                             (iq_ins),
      .valid                           (s2o_valid),
      .op_inv                          (icop_inv),
      .op_inv_paddr                    (icop_inv_paddr),
      .op_stall_req                    (icop_stall_req),
   )
*/
   icache
   #(/*AUTOINSTPARAM*/
     // Parameters
     .CONFIG_AW                         (CONFIG_AW),
     .CONFIG_P_FETCH_WIDTH              (CONFIG_P_FETCH_WIDTH),
     .CONFIG_P_PAGE_SIZE                (CONFIG_P_PAGE_SIZE),
     .CONFIG_IC_P_LINE                  (CONFIG_IC_P_LINE),
     .CONFIG_IC_P_SETS                  (CONFIG_IC_P_SETS),
     .CONFIG_IC_P_WAYS                  (CONFIG_IC_P_WAYS),
     .AXI_P_DW_BYTES                    (AXI_P_DW_BYTES),
     .AXI_ADDR_WIDTH                    (AXI_ADDR_WIDTH),
     .AXI_ID_WIDTH                      (AXI_ID_WIDTH),
     .AXI_USER_WIDTH                    (AXI_USER_WIDTH))
   U_ICACHE
   (/*AUTOINST*/
    // Outputs
    .stall_req                          (ic_stall_req),          // Templated
    .op_stall_req                       (icop_stall_req),        // Templated
    .ins                                (iq_ins),                // Templated
    .valid                              (s2o_valid),             // Templated
    .axi_ar_valid_o                     (axi_ar_valid_o),
    .axi_ar_addr_o                      (axi_ar_addr_o[AXI_ADDR_WIDTH-1:0]),
    .axi_ar_prot_o                      (axi_ar_prot_o[2:0]),
    .axi_ar_id_o                        (axi_ar_id_o[AXI_ID_WIDTH-1:0]),
    .axi_ar_user_o                      (axi_ar_user_o[AXI_USER_WIDTH-1:0]),
    .axi_ar_len_o                       (axi_ar_len_o[7:0]),
    .axi_ar_size_o                      (axi_ar_size_o[2:0]),
    .axi_ar_burst_o                     (axi_ar_burst_o[1:0]),
    .axi_ar_lock_o                      (axi_ar_lock_o),
    .axi_ar_cache_o                     (axi_ar_cache_o[3:0]),
    .axi_ar_qos_o                       (axi_ar_qos_o[3:0]),
    .axi_ar_region_o                    (axi_ar_region_o[3:0]),
    .axi_r_ready_o                      (axi_r_ready_o),
    // Inputs
    .clk                                (clk),
    .rst                                (rst),
    .vpo                                (vpo[CONFIG_P_PAGE_SIZE-1:0]),
    .ppn_s2                             (ppn_s2[CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0]),
    .kill_req_s2                        (kill_req_s2),
    .op_inv                             (icop_inv),              // Templated
    .op_inv_paddr                       (icop_inv_paddr),        // Templated
    .axi_ar_ready_i                     (axi_ar_ready_i),
    .axi_r_valid_i                      (axi_r_valid_i),
    .axi_r_data_i                       (axi_r_data_i[(1<<AXI_P_DW_BYTES)*8-1:0]),
    .axi_r_resp_i                       (axi_r_resp_i[1:0]),
    .axi_r_last_i                       (axi_r_last_i),
    .axi_r_id_i                         (axi_r_id_i[AXI_ID_WIDTH-1:0]),
    .axi_r_user_i                       (axi_r_user_i[AXI_USER_WIDTH-1:0]));

   bpu
      #(/*AUTOINSTPARAM*/
        // Parameters
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH))
   U_BPU
      (
         .clk                           (clk),
         .rst                           (rst),
         .re                            (p_ce),
         .pc                            (s1i_bpu_pc),
         .npc                           (s1o_bpu_npc_packed),
         .upd                           (s1o_bpu_upd_packed),
         // WB
         .bpu_wb                        (bpu_wb),
         .bpu_wb_is_bcc                 (bpu_wb_is_bcc),
         .bpu_wb_is_breg                (bpu_wb_is_breg),
         .bpu_wb_bcc_taken              (bpu_wb_bcc_taken),
         .bpu_wb_pc                     (bpu_wb_pc),
         .bpu_wb_npc_act                (bpu_wb_npc_act),
         .bpu_wb_upd                    (bpu_wb_upd)
      );

   // Collect branch predication info
   generate
      for(i=0;i<FW;i=i+1)
         begin
            assign s1i_bpu_pc[i*(CONFIG_AW-2) +: (CONFIG_AW-2)] = s1i_pc[i][CONFIG_AW-1:2]; // Aligned at 4byte boundary
            assign s1o_bpu_upd[i] = s1o_bpu_upd_packed[i*`BPU_UPD_W +: `BPU_UPD_W];
            assign s1o_bpu_taken[i] = s1o_bpu_upd[i][`BPU_UPD_TAKEN];
            assign s1o_bpu_npc[i] = s1o_bpu_npc_packed[i*(CONFIG_AW-2) +: (CONFIG_AW-2)];
         end
   endgenerate

   priority_encoder  #(.P_DW (CONFIG_P_FETCH_WIDTH)) U_ENC_BP (.din(s1o_bpu_taken), .dout(s1o_bpu_taken_inst_idx) );

   // Generate valid mask
   always @(*)
      begin
         s1i_valid_msk[0] = 'b1;
         for(j=1;j<FW;j=j+1)
            s1i_valid_msk[j] = s1i_valid_msk[j-1] & ~s1o_bpu_taken[j-1];
      end
   
   // Process unaligned access
   generate
      for(i=0;i<FW;i=i+1)
         assign s1i_fetch_valid[i] = (pc_nxt[`NCPU_P_INSN_LEN +: CONFIG_P_FETCH_WIDTH] <= i);
   endgenerate
   
   assign pred_branch_taken = (|s1o_bpu_taken);
   
   // NPC Generator
   always @(*)
      if (flush)
         pc_nxt = flush_tgt;
      else if (~p_ce)
         pc_nxt = pc;
      else if (pred_branch_taken)
         pc_nxt = {s1o_bpu_npc[s1o_bpu_taken_inst_idx], 2'b00};
      else
         pc_nxt = pc + {{CONFIG_AW-CONFIG_P_FETCH_WIDTH-1-`NCPU_P_INSN_LEN{1'b0}}, s1o_push_cnt, {`NCPU_P_INSN_LEN{1'b0}}};

   // PC Register
   mDFF_r # (.DW(CONFIG_AW)) ff_pc (.CLK(clk), .RST(rst), .D(pc_nxt), .Q(pc) );

   assign p_ce = (~ic_stall_req & iq_ready);
   
   assign s1i_fetch_vaddr = {pc_nxt[CONFIG_AW-1:P_FETCH_DW_BYTES], {P_FETCH_DW_BYTES{1'b0}}}; // Aligned by fetch window
   
   // Count the number of valid inst
   clo #(.P_DW(CONFIG_P_FETCH_WIDTH)) U_CLO (.bitmap(s1i_fetch_valid & s1i_valid_msk), .count(s1i_push_cnt) );
   
   assign vpo = s1i_fetch_vaddr[CONFIG_P_PAGE_SIZE-1:0];
   
   // TODO: TLB
   mDFF_r # (.DW(CONFIG_AW-CONFIG_P_PAGE_SIZE)) ff_ppn_s2 (.CLK(clk), .RST(rst), .D(s1i_fetch_vaddr[CONFIG_P_PAGE_SIZE +: CONFIG_AW-CONFIG_P_PAGE_SIZE]), .Q(ppn_s2) );
   assign kill_req_s2 = 'b0;
   assign s1o_exc = 'b0;

   // Control path
   mDFF_lr # (.DW(CONFIG_P_FETCH_WIDTH+1)) ff_s1o_push_cnt (.CLK(clk), .RST(rst), .LOAD(p_ce|flush), .D(s1i_push_cnt & {CONFIG_P_FETCH_WIDTH+1{~flush}}), .Q(s1o_push_cnt) );
   mDFF_lr # (.DW(CONFIG_P_FETCH_WIDTH+1)) ff_s2o_push_cnt (.CLK(clk), .RST(rst), .LOAD(p_ce|flush), .D(s1o_push_cnt & {CONFIG_P_FETCH_WIDTH+1{~flush}}), .Q(s2o_push_cnt) );
   
   // Data path
   mDFF_lr # (.DW(`FNT_EXC_W)) ff_s2o_exc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_exc), .Q(s2o_exc) );
   
   generate
      for(i=0;i<FW;i=i+1)
         begin
            assign s1i_pc[i] = pc_nxt + (i<<`NCPU_P_INSN_LEN);
         
            mDFF_lr # (.DW(CONFIG_AW)) ff_s1o_pc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1i_pc[i]), .Q(s1o_pc[i]) );
            mDFF_lr # (.DW(CONFIG_AW)) ff_s2o_pc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_pc[i]), .Q(s2o_pc[i]) );
            mDFF_lr # (.DW(`BPU_UPD_W)) ff_s2o_bpu_upd (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_bpu_upd[i]), .Q(s2o_bpu_upd[i]) );
            
            assign iq_pc[i*CONFIG_AW +: CONFIG_AW] = s2o_pc[i];
            assign iq_exc[i*`FNT_EXC_W +: `FNT_EXC_W] = s2o_exc;
            assign iq_bpu_upd[i*`BPU_UPD_W +: `BPU_UPD_W] = s2o_bpu_upd[i];
         end
   endgenerate
   
   assign iq_push_cnt = (s2o_push_cnt & {CONFIG_P_FETCH_WIDTH+1{s2o_valid & p_ce}});
   
   // Fetch Buffer
   iq
   #(/*AUTOINSTPARAM*/
     // Parameters
     .CONFIG_AW                         (CONFIG_AW),
     .CONFIG_P_FETCH_WIDTH              (CONFIG_P_FETCH_WIDTH),
     .CONFIG_P_ISSUE_WIDTH              (CONFIG_P_ISSUE_WIDTH),
     .CONFIG_P_IQ_DEPTH                 (CONFIG_P_IQ_DEPTH),
     .CONFIG_PHT_P_NUM                  (CONFIG_PHT_P_NUM),
     .CONFIG_BTB_P_NUM                  (CONFIG_BTB_P_NUM))
   U_IQ
   (/*AUTOINST*/
    // Outputs
    .iq_ready                           (iq_ready),
    .id_valid                           (id_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
    .id_ins                             (id_ins[`NCPU_INSN_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
    .id_pc                              (id_pc[CONFIG_AW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
    .id_exc                             (id_exc[`FNT_EXC_W*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
    .id_bpu_upd                         (id_bpu_upd[`BPU_UPD_W*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
    // Inputs
    .clk                                (clk),
    .rst                                (rst),
    .flush                              (flush),
    .iq_ins                             (iq_ins[`NCPU_INSN_DW*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
    .iq_pc                              (iq_pc[CONFIG_AW*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
    .iq_exc                             (iq_exc[`FNT_EXC_W*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
    .iq_bpu_upd                         (iq_bpu_upd[`BPU_UPD_W*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
    .iq_push_cnt                        (iq_push_cnt[CONFIG_P_FETCH_WIDTH:0]),
    .id_pop_cnt                         (id_pop_cnt[CONFIG_P_ISSUE_WIDTH:0]));
   
endmodule
