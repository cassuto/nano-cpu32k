import "DPI-C" function void dpic_regfile(
   input int r0,
   input int r1,
   input int r2,
   input int r3,
   input int r4,
   input int r5,
   input int r6,
   input int r7,
   input int r8,
   input int r9,
   input int r10,
   input int r11,
   input int r12,
   input int r13,
   input int r14,
   input int r15,
   input int r16,
   input int r17,
   input int r18,
   input int r19,
   input int r20,
   input int r21,
   input int r22,
   input int r23,
   input int r24,
   input int r25,
   input int r26,
   input int r27,
   input int r28,
   input int r29,
   input int r30,
   input int r31
);

module difftest_regfile
(
   input clk,
   input [31:0] r0,
   input [31:0] r1,
   input [31:0] r2,
   input [31:0] r3,
   input [31:0] r4,
   input [31:0] r5,
   input [31:0] r6,
   input [31:0] r7,
   input [31:0] r8,
   input [31:0] r9,
   input [31:0] r10,
   input [31:0] r11,
   input [31:0] r12,
   input [31:0] r13,
   input [31:0] r14,
   input [31:0] r15,
   input [31:0] r16,
   input [31:0] r17,
   input [31:0] r18,
   input [31:0] r19,
   input [31:0] r20,
   input [31:0] r21,
   input [31:0] r22,
   input [31:0] r23,
   input [31:0] r24,
   input [31:0] r25,
   input [31:0] r26,
   input [31:0] r27,
   input [31:0] r28,
   input [31:0] r29,
   input [31:0] r30,
   input [31:0] r31
);

   always @(posedge clk)
      dpic_regfile(
         r0,
         r1,
         r2,
         r3,
         r4,
         r5,
         r6,
         r7,
         r8,
         r9,
         r10,
         r11,
         r12,
         r13,
         r14,
         r15,
         r16,
         r17,
         r18,
         r19,
         r20,
         r21,
         r22,
         r23,
         r24,
         r25,
         r26,
         r27,
         r28,
         r29,
         r30,
         r31
      );

endmodule

