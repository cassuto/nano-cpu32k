library verilog;
use verilog.vl_types.all;
entity tb_ncpu32k_sram is
end tb_ncpu32k_sram;
