// Generator : scripts/build.py
// Toplevel : ysyx_20210479
// Prefix : ysyx_20210479_
// Git hash  : 3dce1fed08158109ac1af930b24e61509ccfa549

module ysyx_20210479_bpu
#(
   parameter                                    CONFIG_PHT_P_NUM = 0,
   parameter                                    CONFIG_BTB_P_NUM = 0,
   parameter                                    CONFIG_AW = 0,
   parameter                                    CONFIG_P_FETCH_WIDTH = 0
)
(
   input                                        clk,
   input                                        rst,
   input                                        re,
   input [(1<<CONFIG_P_FETCH_WIDTH)-1:0]        valid,
   input [(CONFIG_AW-2 )*(1<<CONFIG_P_FETCH_WIDTH)-1:0]  pc,
   output [(CONFIG_AW-2 )*(1<<CONFIG_P_FETCH_WIDTH)-1:0] npc,
   output [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_FETCH_WIDTH)-1:0] upd,
   input                                        bpu_wb,
   input                                        bpu_wb_is_bcc,
   input                                        bpu_wb_is_breg,
   input                                        bpu_wb_is_brel,
   input                                        bpu_wb_taken,
   input [(CONFIG_AW-2 )-1:0]                            bpu_wb_pc,
   input [(CONFIG_AW-2 )-1:0]                            bpu_wb_npc_act,
   input [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]                       bpu_wb_upd
);
   localparam PHT_NUM                           = (1<<CONFIG_PHT_P_NUM);
   localparam BTB_NUM                           = (1<<CONFIG_BTB_P_NUM);
   localparam PHT_DW                            = 2; 
   localparam BTB_DW                            = (1 + 1 + CONFIG_AW-CONFIG_BTB_P_NUM-2 + (CONFIG_AW-2 )); 
   wire [(CONFIG_AW-2 )-1:0]                             s1i_pc         [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [(1<<CONFIG_P_FETCH_WIDTH)*CONFIG_PHT_P_NUM-1:0] s1i_pht_addr;
   wire [(1<<CONFIG_P_FETCH_WIDTH)*CONFIG_BTB_P_NUM-1:0] s1i_btb_addr;
   wire [(CONFIG_AW-2 )-1:0]                             s1o_pc         [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [CONFIG_PHT_P_NUM-1:0]                  s1o_pht_addr   [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [CONFIG_BTB_P_NUM-1:0]                  s1o_btb_addr   [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [(1<<CONFIG_P_FETCH_WIDTH)*PHT_DW-1:0]  s1o_pht_count;
   wire [PHT_DW-1:0]                            s2i_pht_count  [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire                                         s2i_pht_taken  [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [(1<<CONFIG_P_FETCH_WIDTH)*BTB_DW-1:0]  s1o_btb_data;
   wire                                         s2i_btb_v      [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire                                         s2i_btb_is_bcc [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [CONFIG_AW-CONFIG_BTB_P_NUM-3:0]        s2i_btb_tag    [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [(CONFIG_AW-2 )-1:0]                             s2i_btb_npc    [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire                                         s2i_btb_hit    [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire                                         s2i_taken      [(1<<CONFIG_P_FETCH_WIDTH)-1:0];
   wire [CONFIG_PHT_P_NUM-1:0]                  wb_pht_addr;
   wire [CONFIG_BTB_P_NUM-1:0]                  wb_btb_addr;
   wire [PHT_DW-1:0]                            wb_pht_count_org;
   wire                                         wb_pht_we;
   reg [PHT_DW-1:0]                             wb_pht_din;
   wire                                         wb_btb_we;
   wire [BTB_DW-1:0]                            wb_btb_din;
   wire                                         wb_pred_taken; 
   wire [(CONFIG_AW-2 )-1:0]                             wb_pred_tgt; 
   wire [CONFIG_PHT_P_NUM-1:0]                  GHSR_ff;
   wire [CONFIG_PHT_P_NUM-1:0]                  GHSR_nxt;
   genvar i;
   generate
      for(i=0;i<(1<<CONFIG_P_FETCH_WIDTH);i=i+1)
         begin
            ysyx_20210479_mDFF_l #(.DW((CONFIG_AW-2 ))) ff_s1o_pc (.CLK(clk), .LOAD(re), .D(s1i_pc[i]), .Q(s1o_pc[i]) );
            ysyx_20210479_mDFF_l #(.DW(CONFIG_PHT_P_NUM)) ff_s1o_pht_addr (.CLK(clk), .LOAD(re), .D(s1i_pht_addr[i*CONFIG_PHT_P_NUM +: CONFIG_PHT_P_NUM]), .Q(s1o_pht_addr[i]) );
            ysyx_20210479_mDFF_l #(.DW(CONFIG_BTB_P_NUM)) ff_s1o_btb_addr (.CLK(clk), .LOAD(re), .D(s1i_btb_addr[i*CONFIG_BTB_P_NUM +: CONFIG_BTB_P_NUM]), .Q(s1o_btb_addr[i]) );
            assign s1i_pc[i] = pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )];
            assign s1i_pht_addr[i*CONFIG_PHT_P_NUM +: CONFIG_PHT_P_NUM] = s1i_pc[i][CONFIG_PHT_P_NUM-1:0] ^ GHSR_ff;
            assign s1i_btb_addr[i*CONFIG_BTB_P_NUM +: CONFIG_BTB_P_NUM] = s1i_pc[i][CONFIG_BTB_P_NUM-1:0];
            assign s2i_pht_count[i] = s1o_pht_count[i*PHT_DW +: PHT_DW];
            assign s2i_pht_taken[i] = s2i_pht_count[i][PHT_DW-1];
            assign {s2i_btb_npc[i], s2i_btb_tag[i], s2i_btb_is_bcc[i], s2i_btb_v[i]} = s1o_btb_data[i*BTB_DW +: BTB_DW];
            assign s2i_btb_hit[i] = (s2i_btb_v[i] & (s2i_btb_tag[i] == s1o_pc[i][(CONFIG_AW-2 )-1:CONFIG_BTB_P_NUM]));
            assign s2i_taken[i] = (valid[i] & (s2i_btb_hit[i] & (~s2i_btb_is_bcc[i] | s2i_pht_taken[i])));
            assign npc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )] = s2i_btb_npc[i];
            assign upd[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)] = {s1o_pht_count[i*PHT_DW +: PHT_DW], s1o_pht_addr[i], s1o_btb_addr[i], s2i_btb_npc[i], s2i_taken[i]};
         end
   endgenerate
   ysyx_20210479_mRF_nwnr
      #(
         .DW         (PHT_DW),
         .AW         (CONFIG_PHT_P_NUM),
         .NUM_READ   (1<<CONFIG_P_FETCH_WIDTH),
         .NUM_WRITE  (1)
      )
   U_PHT
      (
         .CLK        (clk),
         .RE         ({(1<<CONFIG_P_FETCH_WIDTH){re}}),
         .RADDR      (s1i_pht_addr),
         .RDATA      (s1o_pht_count),
         .WE         (wb_btb_we),
         .WADDR      (wb_pht_addr),
         .WDATA      (wb_pht_din)
      );
   ysyx_20210479_mRF_nwnr
      #(
         .DW         (BTB_DW),
         .AW         (CONFIG_BTB_P_NUM),
         .NUM_READ   (1<<CONFIG_P_FETCH_WIDTH),
         .NUM_WRITE  (1)
      )
   U_BTB
      (
         .CLK        (clk),
         .RE         ({((1<<CONFIG_P_FETCH_WIDTH)){re}}),
         .RADDR      (s1i_btb_addr),
         .RDATA      (s1o_btb_data),
         .WE         (wb_btb_we),
         .WADDR      (wb_btb_addr),
         .WDATA      (wb_btb_din)
      );
   assign {wb_pht_count_org, wb_pht_addr, wb_btb_addr, wb_pred_tgt, wb_pred_taken} = bpu_wb_upd;
   assign wb_pht_we = (bpu_wb & bpu_wb_is_bcc);
   always @(*)
      if (bpu_wb_taken)
         wb_pht_din = (wb_pht_count_org == 2'b11)
                        ? 2'b11
                        : wb_pht_count_org + 'b1;
      else
         wb_pht_din =  (wb_pht_count_org == 2'b00)
                        ? 2'b00
                        : wb_pht_count_org - 'b1;
   assign wb_btb_we = (bpu_wb & (bpu_wb_is_breg | bpu_wb_is_brel));
   assign wb_btb_din = {bpu_wb_npc_act, bpu_wb_pc[(CONFIG_AW-2 )-1:CONFIG_BTB_P_NUM], bpu_wb_is_bcc, 1'b1};
   assign GHSR_nxt = wb_pht_we ? {GHSR_ff[CONFIG_PHT_P_NUM-2:0], bpu_wb_taken}: GHSR_ff;
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_PHT_P_NUM)) ff_GHSR (.CLK(clk), .RST(rst), .LOAD(wb_pht_we), .D(GHSR_nxt), .Q(GHSR_ff) );
endmodule
module ysyx_20210479_cmt
#(
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_ISSUE_WIDTH = 0
)
(
   input                               clk,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_wdat,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_waddr,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)*2-1:0] arf_RE,
   input [(1<<CONFIG_P_ISSUE_WIDTH)*2*5-1:0] arf_RADDR,
   output [(1<<CONFIG_P_ISSUE_WIDTH)*2*CONFIG_DW-1:0] arf_RDATA
);
   localparam IW                       = (1<<CONFIG_P_ISSUE_WIDTH);
   ysyx_20210479_mRF_nwnr
      #(
         .DW                           (CONFIG_DW),
         .AW                           (5),
         .NUM_READ                     (2*IW), 
         .NUM_WRITE                    (IW)
      )
   U_ARF
      (
         .CLK                          (clk),
         .RE                           (arf_RE),
         .RADDR                        (arf_RADDR),
         .RDATA                        (arf_RDATA),
         .WE                           (commit_rf_we),
         .WADDR                        (commit_rf_waddr),
         .WDATA                        (commit_rf_wdat)
      );
endmodule
module ysyx_20210479_dcache
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_DW = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_DC_P_LINE = 0,
   parameter                           CONFIG_DC_P_SETS = 0,
   parameter                           CONFIG_DC_P_WAYS = 0,
   parameter                           AXI_P_DW_BYTES    = 0,
   parameter                           AXI_ADDR_WIDTH    = 0,
   parameter                           AXI_ID_WIDTH      = 0,
   parameter                           AXI_USER_WIDTH    = 0
)
(
   input                               clk,
   input                               rst,
   output                              stall_req,
   input                               req,
   input [2:0]                         size,
   input [CONFIG_DW/8-1:0]             wmsk,
   input [CONFIG_DW-1:0]               wdat,
   input [CONFIG_P_PAGE_SIZE-1:0]      vpo,
   input [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] ppn_s2,
   input                               kill_req_s2,
   input                               uncached_s2,
   input                               inv,
   input                               fls,
   output [CONFIG_DW-1:0]              dout,
   input                               dbus_ARREADY,
   output                              dbus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_ARADDR,
   output [2:0]                        dbus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_ARID,
   output [AXI_USER_WIDTH-1:0]         dbus_ARUSER,
   output [7:0]                        dbus_ARLEN,
   output [2:0]                        dbus_ARSIZE,
   output [1:0]                        dbus_ARBURST,
   output                              dbus_ARLOCK,
   output [3:0]                        dbus_ARCACHE,
   output [3:0]                        dbus_ARQOS,
   output [3:0]                        dbus_ARREGION,
   output                              dbus_RREADY,
   input                               dbus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_RDATA,
   input                               dbus_RLAST,
   input                               dbus_AWREADY,
   output                              dbus_AWVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_AWADDR,
   output [2:0]                        dbus_AWPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_AWID,
   output [AXI_USER_WIDTH-1:0]         dbus_AWUSER,
   output [7:0]                        dbus_AWLEN,
   output [2:0]                        dbus_AWSIZE,
   output [1:0]                        dbus_AWBURST,
   output                              dbus_AWLOCK,
   output [3:0]                        dbus_AWCACHE,
   output [3:0]                        dbus_AWQOS,
   output [3:0]                        dbus_AWREGION,
   input                               dbus_WREADY,
   output                              dbus_WVALID,
   output [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_WDATA,
   output [(1<<AXI_P_DW_BYTES)-1:0]    dbus_WSTRB,
   output                              dbus_WLAST,
   output [AXI_USER_WIDTH-1:0]         dbus_WUSER,
   output                              dbus_BREADY,
   input                               dbus_BVALID,
   input  [1:0]                        dbus_RRESP, 
   input  [AXI_ID_WIDTH-1:0]           dbus_RID, 
   input  [AXI_USER_WIDTH-1:0]         dbus_RUSER, 
   input [1:0]                         dbus_BRESP, 
   input [AXI_ID_WIDTH-1:0]            dbus_BID, 
   input [AXI_USER_WIDTH-1:0]          dbus_BUSER, 
   output [CONFIG_DW-1:0]              msr_dcid
);
   localparam TAG_WIDTH                = (CONFIG_AW - CONFIG_DC_P_SETS - CONFIG_DC_P_LINE);
   localparam TAG_V_RAM_AW             = (CONFIG_DC_P_SETS);
   localparam TAG_V_RAM_DW             = (TAG_WIDTH + 1); 
   localparam PAYLOAD_DW               = (CONFIG_DW);
   localparam PAYLOAD_P_DW_BYTES       = (CONFIG_P_DW-3); 
   localparam PAYLOAD_AW               = (CONFIG_DC_P_SETS + CONFIG_DC_P_LINE - PAYLOAD_P_DW_BYTES);
   localparam AXI_FETCH_SIZE           = (PAYLOAD_P_DW_BYTES <= AXI_P_DW_BYTES) ? PAYLOAD_P_DW_BYTES : AXI_P_DW_BYTES;
   reg [CONFIG_DC_P_SETS-1:0]          s1i_line_addr;
   reg [TAG_V_RAM_DW-1:0]              s1i_replace_tag_v;
   wire                                s1i_tag_v_re;
   wire                                s1i_tag_v_we            [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire                                s1o_inv;
   wire                                s1o_fls;
   reg                                 s2i_ready;
   wire                                s2i_d_we                [(1<<CONFIG_DC_P_WAYS)-1:0];
   reg [TAG_V_RAM_AW-1:0]              s2i_d_waddr;
   reg                                 s2i_d_wdat              [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire [PAYLOAD_DW/8-1:0]             s2i_payload_we          [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire [PAYLOAD_DW/8-1:0]             s2i_payload_tgt_we;
   reg [PAYLOAD_DW-1:0]                s2i_payload_din;
   wire [PAYLOAD_DW/8-1:0]             s2i_wb_we;
   wire [PAYLOAD_DW-1:0]               s2i_wb_din;
   wire                                s2i_wb_re;
   wire [2:0]                          s1o_size;
   wire [CONFIG_DW/8-1:0]              s1o_wmsk;
   wire [CONFIG_DW-1:0]                s1o_wdat;
   wire [CONFIG_DC_P_SETS-1:0]         s1o_line_addr;
   reg [PAYLOAD_AW-1:0]                s2i_payload_addr;
   wire                                s2i_payload_re;
   wire                                s1o_valid;
   wire [TAG_V_RAM_DW-1:0]             s1o_tag_v               [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s1o_d;
   wire                                s1o_free_dirty;
   wire [TAG_WIDTH-1:0]                s2i_free_tag;
   wire [CONFIG_P_PAGE_SIZE-1:0]       s1o_vpo;
   wire [CONFIG_AW-1:0]                s2i_paddr;
   wire [TAG_WIDTH-1:0]                s2i_tag                 [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire [TAG_WIDTH*(1<<CONFIG_DC_P_WAYS)-1:0] s2i_tag_packed;
   wire                                s2i_v                   [(1<<CONFIG_DC_P_WAYS)-1:0];
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2i_hit_vec;
   wire                                s2i_hit;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2i_match_vec;
   wire                                s2i_match_vec_ce;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2o_fsm_free_way;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2i_wb_way;
   wire                                s2o_fls;
   wire [CONFIG_DC_P_SETS-1:0]         s2o_line_addr;
   wire [CONFIG_AW-1:0]                s2o_paddr;
   wire [CONFIG_DW/8-1:0]              s2o_wmsk;
   wire [CONFIG_DW-1:0]                s2o_wdat;
   wire [PAYLOAD_DW*(1<<CONFIG_DC_P_WAYS)-1:0] s2o_payload;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2o_match_vec;
   wire [PAYLOAD_DW-1:0]               s2o_match_payload;
   wire [PAYLOAD_DW-1:0]               s2o_wb_payload;
   wire                                s2o_free_dirty;
   wire [TAG_WIDTH-1:0]                s2o_free_tag;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    s2o_d;
   wire                                s2o_match_dirty;
   wire [PAYLOAD_AW-1:0]               s2o_payload_addr;
   wire [CONFIG_DC_P_LINE-1:0]         s2o_wb_addr;
   wire [2:0]                          s2o_size;
   wire                                s2o_uncached;
   reg [3:0]                           fsm_state_nxt;
   wire [3:0]                          fsm_state_ff;
   wire [(1<<CONFIG_DC_P_WAYS)-1:0]    fsm_free_way, fsm_free_way_nxt;
   wire [CONFIG_DC_P_SETS-1:0]         fsm_boot_cnt;
   wire [CONFIG_DC_P_SETS:0]           fsm_boot_cnt_nxt_carry;
   wire [CONFIG_DC_P_LINE-1:0]         fsm_refill_cnt;
   wire [CONFIG_DC_P_LINE:0]           fsm_refill_cnt_nxt_carry;
   reg [CONFIG_DC_P_LINE-1:0]          fsm_refill_cnt_nxt;
   reg                                 fsm_uncached_req;
   wire                                p_ce;
   wire [CONFIG_AW-1:0]                axi_paddr_nxt;
   reg                                 ar_set, aw_set;
   wire                                ar_clr, aw_clr;
   wire                                wvalid_set, wvalid_clr;
   wire                                wlast_set, wlast_clr;
   wire                                hds_axi_R;
   wire                                hds_axi_R_last;
   wire                                hds_axi_W;
   wire                                hds_axi_W_last;
   wire                                hds_axi_B;
   wire [AXI_ADDR_WIDTH-1:0]           axi_arw_addr_nxt;
   wire [PAYLOAD_DW-1:0]               axi_aligned_rdata_ff;
   wire [PAYLOAD_DW/8-1:0]             axi_aligned_rdata_ff_wmsk;
   wire [PAYLOAD_DW-1:0]               axi_aligned_rdata_nxt;
   localparam [3:0] S_BOOT             = 4'd0;
   localparam [3:0] S_IDLE             = 4'd1;
   localparam [3:0] S_REPLACE          = 4'd2;
   localparam [3:0] S_REFILL           = 4'd3;
   localparam [3:0] S_WRITEBACK        = 4'd4;
   localparam [3:0] S_INVALIDATE       = 4'd5;
   localparam [3:0] S_RELOAD_S1O_S2O   = 4'd6;
   localparam [3:0] S_FLUSH            = 4'd7;
   localparam [3:0] S_UNCACHED_BOOT    = 4'd8;
   localparam [3:0] S_UNCACHED_READ    = 4'd9;
   localparam [3:0] S_UNCACHED_WRITE   = 4'd10;
   genvar way, i, j;
   assign p_ce = (~stall_req);
   generate
      for(way=0; way<(1<<CONFIG_DC_P_WAYS); way=way+1)
         begin : gen_ways
            wire rf_d, rf_d_ff;
            wire rf_conflict;
            wire rf_bypass;
            ysyx_20210479_mRAM_s_s_be
               #(
                  .P_DW (PAYLOAD_P_DW_BYTES + 3),
                  .AW   (PAYLOAD_AW)
               )
            U_PAYLOAD_RAM
               (
                  .CLK  (clk),
                  .ADDR (s2i_payload_addr),
                  .RE   (s2i_payload_re),
                  .DOUT (s2o_payload[way*PAYLOAD_DW +: PAYLOAD_DW]),
                  .WE   (s2i_payload_we[way]),
                  .DIN  (s2i_payload_din)
               );
            ysyx_20210479_mRF_1wr
               #(
                  .DW   (TAG_V_RAM_DW),
                  .AW   (TAG_V_RAM_AW)
               )
            U_TAG_V_RAM
               (
                  .CLK  (clk),
                  .ADDR (s1i_line_addr),
                  .RE   (s1i_tag_v_re),
                  .RDATA (s1o_tag_v[way]),
                  .WE   (s1i_tag_v_we[way]),
                  .WDATA (s1i_replace_tag_v)
               );
            ysyx_20210479_mRF_nwnr
               #(
                  .DW   (1),
                  .AW   (TAG_V_RAM_AW),
                  .NUM_READ (1),
                  .NUM_WRITE (1)
               )
            U_D_RF
               (
                  .CLK     (clk),
                  .RE      (s1i_tag_v_re),
                  .RADDR   (s1i_line_addr),
                  .RDATA   (rf_d),
                  .WE      (s2i_d_we[way]),
                  .WADDR   (s2i_d_waddr),
                  .WDATA   (s2i_d_wdat[way])
               );
            assign rf_conflict = ((s1i_line_addr == s2i_d_waddr) & s2i_d_we[way]);
            ysyx_20210479_mDFF_lr #(.DW(1)) ff_bypass (.CLK(clk), .RST(rst), .LOAD(rf_conflict | s1i_tag_v_re), .D(rf_conflict | ~s1i_tag_v_re), .Q(rf_bypass) );
            ysyx_20210479_mDFF_l #(.DW(1)) ff_rd_d (.CLK(clk), .LOAD(s1i_tag_v_re), .D(s2i_d_wdat[way]), .Q(rf_d_ff) );
            assign s1o_d[way] = rf_bypass ? rf_d_ff : rf_d;
            assign {s2i_tag[way], s2i_v[way]} = s1o_tag_v[way];
            assign s2i_tag_packed[way * TAG_WIDTH +: TAG_WIDTH] = s2i_tag[way];
            assign s2i_hit_vec[way] = (s2i_v[way] & (s2i_tag[way] == s2i_paddr[CONFIG_AW-1:CONFIG_DC_P_LINE+CONFIG_DC_P_SETS]) );
         end
   endgenerate
   assign s2i_hit = (|s2i_hit_vec);
   assign s2i_match_vec = (fsm_state_ff==S_RELOAD_S1O_S2O) ? s2o_fsm_free_way : s2i_hit_vec;
   assign s2i_match_vec_ce = (p_ce | (fsm_state_ff==S_RELOAD_S1O_S2O));
   assign s2i_wb_way = (s2o_fls) ? s2o_match_vec : s2o_fsm_free_way;
   ysyx_20210479_pmux #(.SELW(1<<CONFIG_DC_P_WAYS), .DW(PAYLOAD_DW)) pmux_s2o_payload (.sel(s2o_match_vec), .din(s2o_payload), .dout(s2o_match_payload));
   ysyx_20210479_pmux #(.SELW(1<<CONFIG_DC_P_WAYS), .DW(1)) pmux_s2o_d (.sel(s2o_match_vec), .din(s2o_d), .dout(s2o_match_dirty));
   ysyx_20210479_pmux #(.SELW(1<<CONFIG_DC_P_WAYS), .DW(PAYLOAD_DW)) pmux_s2o_wb_payload (.sel(s2i_wb_way), .din(s2o_payload), .dout(s2o_wb_payload));
   ysyx_20210479_pmux #(.SELW(1<<CONFIG_DC_P_WAYS), .DW(1)) pmux_s1o_free_dirty (.sel(fsm_free_way), .din(s1o_d), .dout(s1o_free_dirty));
   ysyx_20210479_pmux #(.SELW(1<<CONFIG_DC_P_WAYS), .DW(TAG_WIDTH)) pmux_s2i_free_tag (.sel(fsm_free_way), .din(s2i_tag_packed), .dout(s2i_free_tag));
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_valid (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(req), .Q(s1o_valid) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_inv (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(inv), .Q(s1o_inv) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_fls (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(fls), .Q(s1o_fls) );
   ysyx_20210479_mDFF_l # (.DW(3)) ff_s1o_size (.CLK(clk), .LOAD(p_ce), .D(size), .Q(s1o_size) );
   ysyx_20210479_mDFF_lr # (.DW(CONFIG_DW/8)) ff_s1o_wmsk (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(wmsk), .Q(s1o_wmsk) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW)) ff_s1o_wdat (.CLK(clk), .LOAD(p_ce), .D(wdat), .Q(s1o_wdat) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_P_PAGE_SIZE)) ff_s1o_vpo (.CLK(clk), .LOAD(p_ce), .D(vpo), .Q(s1o_vpo) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DC_P_SETS)) ff_s1o_line_addr (.CLK(clk), .LOAD(p_ce), .D(s1i_line_addr), .Q(s1o_line_addr) );
   ysyx_20210479_mDFF_l # (.DW(1<<CONFIG_DC_P_WAYS)) ff_s2o_match_vec (.CLK(clk), .LOAD(s2i_match_vec_ce), .D(s2i_match_vec), .Q(s2o_match_vec) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DC_P_SETS)) ff_s2o_line_addr (.CLK(clk), .LOAD(p_ce), .D(s1o_line_addr), .Q(s2o_line_addr) );
   ysyx_20210479_mDFF_l # (.DW(1<<CONFIG_DC_P_WAYS)) ff_s2o_fsm_free_way (.CLK(clk), .LOAD(p_ce), .D(fsm_free_way), .Q(s2o_fsm_free_way) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s2o_fls (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_fls), .Q(s2o_fls) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_AW)) ff_s2o_paddr (.CLK(clk), .LOAD(p_ce), .D(s2i_paddr), .Q(s2o_paddr) );
   ysyx_20210479_mDFF_l # (.DW(1<<CONFIG_DC_P_WAYS)) ff_s2o_d (.CLK(clk), .LOAD(p_ce), .D(s1o_d), .Q(s2o_d) );
   ysyx_20210479_mDFF_l # (.DW(1)) ff_s2o_free_dirty (.CLK(clk), .LOAD(p_ce), .D(s1o_free_dirty), .Q(s2o_free_dirty) );
   ysyx_20210479_mDFF_l # (.DW(TAG_WIDTH)) ff_s2o_free_tag (.CLK(clk), .LOAD(p_ce), .D(s2i_free_tag), .Q(s2o_free_tag) );
   ysyx_20210479_mDFF_l # (.DW(PAYLOAD_AW)) ff_s2o_payload_addr (.CLK(clk), .LOAD(p_ce), .D(s2i_payload_addr), .Q(s2o_payload_addr) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DC_P_LINE)) ff_s2o_wb_addr (.CLK(clk), .LOAD(s2i_wb_re), .D(fsm_refill_cnt), .Q(s2o_wb_addr) );
   ysyx_20210479_mDFF_l # (.DW(3)) ff_s2o_size (.CLK(clk), .LOAD(p_ce), .D(s1o_size), .Q(s2o_size) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW)) ff_s2o_wdat (.CLK(clk), .LOAD(p_ce), .D(s1o_wdat), .Q(s2o_wdat) );
   ysyx_20210479_mDFF_lr # (.DW(CONFIG_DW/8)) ff_s2o_wmsk (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_wmsk), .Q(s2o_wmsk) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s2o_use_uncached_dout (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(uncached_s2), .Q(s2o_uncached) );
   always @(*)
      begin
         fsm_state_nxt = fsm_state_ff;
         ar_set = 'b0;
         aw_set = 'b0;
         fsm_uncached_req = 'b0;
         s2i_ready = 'b0;
         case (fsm_state_ff)
            S_BOOT:
               if (fsm_boot_cnt_nxt_carry[CONFIG_DC_P_SETS])
                  fsm_state_nxt = S_IDLE;
            S_IDLE:
               if (s1o_valid)
                  if (s1o_inv)
                     fsm_state_nxt = S_INVALIDATE;
                  else if (s1o_fls)
                     fsm_state_nxt = s2i_hit ? S_FLUSH : S_IDLE;
                  else if (uncached_s2 & ~kill_req_s2) 
                     fsm_state_nxt = S_UNCACHED_BOOT;
                  else if (~s2i_hit & ~uncached_s2 & ~kill_req_s2) 
                     fsm_state_nxt = S_REPLACE;
                  else if (s2i_hit & ~uncached_s2 & ~kill_req_s2) 
                     s2i_ready = 'b1;
            S_REPLACE:
               begin
                  fsm_state_nxt = (s2o_free_dirty) ? S_WRITEBACK : S_REFILL;
                  ar_set = ~s2o_free_dirty;
                  aw_set = s2o_free_dirty;
               end
            S_WRITEBACK:
               if (hds_axi_B)
                  begin
                     fsm_state_nxt = (s2o_fls) ? S_IDLE : S_REFILL;
                     ar_set = ~s2o_fls;
                  end
            S_REFILL:
               if (hds_axi_R_last)
                  fsm_state_nxt = S_RELOAD_S1O_S2O;
            S_INVALIDATE:
               fsm_state_nxt = S_IDLE;
            S_RELOAD_S1O_S2O:
               fsm_state_nxt = S_IDLE;
            S_FLUSH:
               begin
                  fsm_state_nxt = (s2o_match_dirty) ? S_WRITEBACK : S_IDLE;
                  aw_set = s2o_match_dirty;
               end
            S_UNCACHED_BOOT:
               begin
                  fsm_state_nxt = (|s2o_wmsk) ? S_UNCACHED_WRITE : S_UNCACHED_READ;
                  ar_set = ~(|s2o_wmsk);
                  aw_set = (|s2o_wmsk);
                  fsm_uncached_req = 'b1;
               end
            S_UNCACHED_READ:
               if (hds_axi_R)
                  fsm_state_nxt = S_IDLE;
            S_UNCACHED_WRITE:
               if (hds_axi_B)
                  fsm_state_nxt = S_IDLE;
            default: ;
         endcase
      end
   ysyx_20210479_mDFF_r # (.DW(4), .RST_VECTOR(S_BOOT)) ff_state_r (.CLK(clk), .RST(rst), .D(fsm_state_nxt), .Q(fsm_state_ff) );
   assign fsm_free_way_nxt = (fsm_free_way[(1<<CONFIG_DC_P_WAYS)-1])
                              ? {{(1<<CONFIG_DC_P_WAYS)-1{1'b0}}, 1'b1}
                              : {fsm_free_way[(1<<CONFIG_DC_P_WAYS)-2:0], 1'b0};
   ysyx_20210479_mDFF_r #(.DW(1<<CONFIG_DC_P_WAYS), .RST_VECTOR({{(1<<CONFIG_DC_P_WAYS)-1{1'b0}}, 1'b1}) ) ff_fsm_free_idx
      (.CLK(clk), .RST(rst), .D(fsm_free_way_nxt), .Q(fsm_free_way) );
   assign fsm_boot_cnt_nxt_carry = fsm_boot_cnt + 'b1;
   ysyx_20210479_mDFF_r # (.DW(CONFIG_DC_P_SETS)) ff_fsm_boot_cnt_nxt (.CLK(clk), .RST(rst), .D(fsm_boot_cnt_nxt_carry[CONFIG_DC_P_SETS-1:0]), .Q(fsm_boot_cnt) );
   always @(*)
      if (((fsm_state_ff==S_REFILL) & hds_axi_R) | s2i_wb_re)
         fsm_refill_cnt_nxt = fsm_refill_cnt_nxt_carry[CONFIG_DC_P_LINE-1:0];
      else
         fsm_refill_cnt_nxt = fsm_refill_cnt;
   assign fsm_refill_cnt_nxt_carry = (fsm_refill_cnt + (1<<AXI_FETCH_SIZE));
   ysyx_20210479_mDFF_r # (.DW(CONFIG_DC_P_LINE)) ff_fsm_refill_cnt (.CLK(clk), .RST(rst), .D(fsm_refill_cnt_nxt), .Q(fsm_refill_cnt) );
   always @(*)
      case (fsm_state_ff)
         S_BOOT:
            s1i_line_addr = fsm_boot_cnt;
         S_INVALIDATE,
         S_REPLACE:
            s1i_line_addr = s2o_line_addr;
         S_RELOAD_S1O_S2O:
            s1i_line_addr = s1o_line_addr;
         default:
            s1i_line_addr = vpo[CONFIG_DC_P_LINE +: CONFIG_DC_P_SETS]; 
      endcase
   always @(*)
      case (fsm_state_ff)
         S_REPLACE:
            s1i_replace_tag_v = {s2o_paddr[CONFIG_AW-1:CONFIG_DC_P_LINE+CONFIG_DC_P_SETS], 1'b1};
         default: 
            s1i_replace_tag_v = 'b0;
      endcase
   assign s1i_tag_v_re = (p_ce | (fsm_state_ff==S_RELOAD_S1O_S2O));
   generate
      for(way=0; way<(1<<CONFIG_DC_P_WAYS); way=way+1)
         assign s1i_tag_v_we[way] = (fsm_state_ff==S_BOOT) |
                                    (fsm_state_ff==S_INVALIDATE) |
                                    ((fsm_state_ff==S_REPLACE) & (s2o_fsm_free_way[way]));
   endgenerate
   always @(*)
      case (fsm_state_ff)
         S_IDLE:
            s2i_d_waddr = s1o_line_addr;
         S_RELOAD_S1O_S2O:
            s2i_d_waddr = s2o_line_addr;
         default:
            s2i_d_waddr = s1i_line_addr;
      endcase
   generate
      for(way=0; way<(1<<CONFIG_DC_P_WAYS); way=way+1)
         always @(*)
            case (fsm_state_ff)
               S_IDLE:
                  s2i_d_wdat[way] = s1o_d[way] | (|s1o_wmsk);
               S_RELOAD_S1O_S2O:
                  s2i_d_wdat[way] = s2o_d[way] | (|s2o_wmsk);
               default: 
                  s2i_d_wdat[way] = 'b0;
            endcase
   endgenerate
   generate
      for(way=0; way<(1<<CONFIG_DC_P_WAYS); way=way+1)
         assign s2i_d_we[way] = (fsm_state_ff==S_BOOT) |
                                 (fsm_state_ff==S_INVALIDATE) |
                                 ((fsm_state_ff==S_REPLACE) & (s2o_fsm_free_way[way])) |
                                 ((fsm_state_ff==S_RELOAD_S1O_S2O) & s2o_fsm_free_way[way]) |
                                 (s2i_ready & s2i_hit_vec[way]);
   endgenerate
   assign s2i_paddr = {ppn_s2, s1o_vpo};
   always @(*)
      if (s2i_wb_re)
         s2i_payload_addr = {s2o_paddr[CONFIG_DC_P_LINE +: CONFIG_DC_P_SETS], fsm_refill_cnt[PAYLOAD_P_DW_BYTES +: CONFIG_DC_P_LINE-PAYLOAD_P_DW_BYTES]};
      else
         case (fsm_state_ff)
            S_REFILL:
               s2i_payload_addr = {s2o_paddr[CONFIG_DC_P_LINE +: CONFIG_DC_P_SETS], fsm_refill_cnt[PAYLOAD_P_DW_BYTES +: CONFIG_DC_P_LINE-PAYLOAD_P_DW_BYTES]};
            S_RELOAD_S1O_S2O:
               s2i_payload_addr = s2o_payload_addr;
            default:
               s2i_payload_addr = s1o_vpo[PAYLOAD_P_DW_BYTES +: PAYLOAD_AW]; 
         endcase
   always @(*)
      case (fsm_state_ff)
         S_IDLE:
            s2i_payload_din = s1o_wdat;
         S_RELOAD_S1O_S2O:
            s2i_payload_din = s2o_wdat;
         default:
            s2i_payload_din = s2i_wb_din;
      endcase
   assign s2i_payload_re = (p_ce |
                              s2i_wb_re |
                              (fsm_state_ff==S_RELOAD_S1O_S2O));
   assign s2i_payload_tgt_we = ({CONFIG_DW/8{s2i_ready}} & s1o_wmsk) |
                                 ({CONFIG_DW/8{fsm_state_ff==S_RELOAD_S1O_S2O}} & s2o_wmsk) |
                                 s2i_wb_we;
   generate
      for(way=0;way<(1<<CONFIG_DC_P_WAYS);way=way+1)
         assign s2i_payload_we[way] = (s2i_payload_tgt_we &
                                       {CONFIG_DW/8{
                                          (s2i_ready & s2i_hit_vec[way]) |
                                          ((fsm_state_ff==S_RELOAD_S1O_S2O) & s2o_fsm_free_way[way]) |
                                          ((fsm_state_ff==S_REFILL) & s2o_fsm_free_way[way])
                                       }});
   endgenerate
   ysyx_20210479_align_r
      #(
         .AXI_P_DW_BYTES               (AXI_P_DW_BYTES),
         .PAYLOAD_P_DW_BYTES           (PAYLOAD_P_DW_BYTES),
         .RAM_AW                       (CONFIG_DC_P_LINE)
      )
   U_ALIGN_R
      (
         .i_axi_RDATA                  (dbus_RDATA),
         .i_ram_we                     (fsm_state_ff == S_REFILL),
         .i_ram_addr                   (fsm_refill_cnt),
         .o_ram_wmsk                   (s2i_wb_we),
         .o_ram_din                    (s2i_wb_din)
      );
   assign stall_req = (fsm_state_ff != S_IDLE);
   assign dout = (s2o_uncached)
                     ? axi_aligned_rdata_ff
                     : s2o_match_payload;
   assign dbus_ARPROT = 3'b000 | 3'b000 | 3'b000;
   assign dbus_ARID = {AXI_ID_WIDTH{1'b0}};
   assign dbus_ARUSER = {AXI_USER_WIDTH{1'b0}};
   assign dbus_ARLEN = (fsm_state_ff==S_UNCACHED_READ) ? 'b0 : ((1<<(CONFIG_DC_P_LINE-AXI_FETCH_SIZE))-1);
   assign dbus_ARSIZE = (fsm_state_ff==S_UNCACHED_READ) ? s2o_size : AXI_FETCH_SIZE;
   assign dbus_ARBURST = 2'b01;
   assign dbus_ARLOCK = 'b0;
   assign dbus_ARCACHE = 4'b0010;
   assign dbus_ARQOS = 'b0;
   assign dbus_ARREGION = 'b0;
   assign ar_clr = (dbus_ARREADY & dbus_ARVALID);
   assign axi_paddr_nxt = (fsm_uncached_req)
                           ? 
                              s2o_paddr
                           : ((fsm_state_ff==S_REPLACE) & aw_set)
                              ? 
                                 {s2o_free_tag, s2o_line_addr, {CONFIG_DC_P_LINE{1'b0}}}
                              : 
                                 {s2o_paddr[CONFIG_DC_P_LINE +: CONFIG_AW - CONFIG_DC_P_LINE], {CONFIG_DC_P_LINE{1'b0}}};
   generate
      if (AXI_ADDR_WIDTH > CONFIG_AW)
         assign axi_arw_addr_nxt = {{AXI_ADDR_WIDTH-CONFIG_AW{1'b0}}, axi_paddr_nxt};
      else if (AXI_ADDR_WIDTH < CONFIG_AW)
         assign axi_arw_addr_nxt = axi_paddr_nxt[AXI_ADDR_WIDTH-1:0];
      else
         assign axi_arw_addr_nxt = axi_paddr_nxt;
   endgenerate
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_dbus_ARVALID (.CLK(clk), .RST(rst), .LOAD(ar_set|ar_clr), .D(ar_set|~ar_clr), .Q(dbus_ARVALID) );
   ysyx_20210479_mDFF_lr # (.DW(AXI_ADDR_WIDTH)) ff_dbus_ARADDR (.CLK(clk), .RST(rst), .LOAD(ar_set), .D(axi_arw_addr_nxt), .Q(dbus_ARADDR) );
   assign dbus_RREADY = (fsm_state_ff == S_REFILL) | (fsm_state_ff == S_UNCACHED_READ);
   assign hds_axi_R = (dbus_RVALID & dbus_RREADY);
   assign hds_axi_R_last = (hds_axi_R & dbus_RLAST);
   generate
      if (PAYLOAD_P_DW_BYTES <= AXI_P_DW_BYTES)
         begin : gen_uncached_align
            ysyx_20210479_align_r
               #(
                  .AXI_P_DW_BYTES               (AXI_P_DW_BYTES),
                  .PAYLOAD_P_DW_BYTES           (PAYLOAD_P_DW_BYTES),
                  .RAM_AW                       (AXI_ADDR_WIDTH)
               )
            U_ALIGN_UNUCACHED_R
               (
                  .i_axi_RDATA                  (dbus_RDATA),
                  .i_ram_we                     (hds_axi_R),
                  .i_ram_addr                   (dbus_ARADDR),
                  .o_ram_wmsk                   (axi_aligned_rdata_ff_wmsk),
                  .o_ram_din                    (axi_aligned_rdata_nxt)
               );
            ysyx_20210479_mDFF_l # (.DW(PAYLOAD_DW)) ff_axi_aligned_rdata (.CLK(clk), .LOAD(|axi_aligned_rdata_ff_wmsk), .D(axi_aligned_rdata_nxt), .Q(axi_aligned_rdata_ff) );
         end
      else
         initial $fatal(1, "Unsupported bitwidth for uncached device!");
   endgenerate
   assign dbus_AWPROT = 3'b000 | 3'b000 | 3'b000;
   assign dbus_AWID = {AXI_ID_WIDTH{1'b0}};
   assign dbus_AWUSER = {AXI_USER_WIDTH{1'b0}};
   assign dbus_AWLEN = (fsm_state_ff==S_UNCACHED_WRITE) ? 'b0 : ((1<<(CONFIG_DC_P_LINE-AXI_FETCH_SIZE))-1);
   assign dbus_AWSIZE = (fsm_state_ff==S_UNCACHED_WRITE) ? s2o_size : AXI_FETCH_SIZE;
   assign dbus_AWBURST = 2'b01;
   assign dbus_AWLOCK = 'b0;
   assign dbus_AWCACHE = 4'b0010;
   assign dbus_AWQOS = 'b0;
   assign dbus_AWREGION = 'b0;
   assign aw_clr = (dbus_AWREADY & dbus_AWVALID);
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_dbus_AWVALID (.CLK(clk), .RST(rst), .LOAD(aw_set|aw_clr), .D(aw_set|~aw_clr), .Q(dbus_AWVALID) );
   ysyx_20210479_mDFF_lr # (.DW(AXI_ADDR_WIDTH)) ff_dbus_AWADDR (.CLK(clk), .RST(rst), .LOAD(aw_set), .D(axi_arw_addr_nxt), .Q(dbus_AWADDR) );
   assign dbus_WUSER = 'b0;
   ysyx_20210479_align_w
      #(
         .AXI_P_DW_BYTES                     (AXI_P_DW_BYTES),
         .PAYLOAD_P_DW_BYTES                 (PAYLOAD_P_DW_BYTES),
         .I_AXI_ADDR_AW                      (CONFIG_DC_P_LINE)
      )
   U_ALIGN_W
      (
         .i_axi_din                          ((fsm_state_ff == S_WRITEBACK) ? s2o_wb_payload : s2o_wdat),
         .i_axi_we                           ((fsm_state_ff == S_WRITEBACK) | (fsm_state_ff == S_UNCACHED_WRITE)),
         .i_axi_addr                         ((fsm_state_ff == S_WRITEBACK) ? s2o_wb_addr : dbus_AWADDR[CONFIG_DC_P_LINE-1:0]),
         .o_axi_WSTRB                        (dbus_WSTRB),
         .o_axi_WDATA                        (dbus_WDATA)
      );
   assign s2i_wb_re = (((fsm_state_ff!=S_UNCACHED_BOOT) & wvalid_set) |
                        ((fsm_state_ff==S_WRITEBACK) & hds_axi_W & (|fsm_refill_cnt)));
   assign wvalid_set = (aw_set);
   assign wvalid_clr = (hds_axi_W_last);
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_dbus_WVALID (.CLK(clk), .RST(rst), .LOAD(wvalid_set|wvalid_clr), .D(wvalid_set|~wvalid_clr), .Q(dbus_WVALID) );
   assign wlast_set = (((fsm_state_ff==S_WRITEBACK) & hds_axi_W & fsm_refill_cnt_nxt_carry[CONFIG_DC_P_LINE]) | fsm_uncached_req);
   assign wlast_clr = (wvalid_clr);
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_dbus_WLAST (.CLK(clk), .RST(rst), .LOAD(wlast_set|wlast_clr), .D(wlast_set|~wlast_clr), .Q(dbus_WLAST) );
   assign hds_axi_W = (dbus_WVALID & dbus_WREADY);
   assign hds_axi_W_last = (hds_axi_W & dbus_WLAST);
   assign dbus_BREADY = (fsm_state_ff == S_WRITEBACK) | (fsm_state_ff == S_UNCACHED_WRITE);
   assign hds_axi_B = (dbus_BREADY & dbus_BVALID);
   assign msr_dcid[3:0] = CONFIG_DC_P_SETS[3:0];
   assign msr_dcid[7:4] = CONFIG_DC_P_LINE[3:0];
   assign msr_dcid[11:8] = CONFIG_DC_P_WAYS[3:0];
   assign msr_dcid[31:12] = 20'b0;
endmodule
module ysyx_20210479_dmmu
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_DMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_DTLB_P_SETS = 0
)
(
   input                               clk,
   input                               rst,
   input                               re,
   input [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] vpn,
   input                               we,
   output [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] ppn,
   output                              EDTM,
   output                              EDPF,
   output                              uncached,
   input                               msr_psr_dmme,
   input                               msr_psr_rm,
   output [CONFIG_DW-1:0]              msr_dmmid,
   input [CONFIG_DTLB_P_SETS-1:0]      msr_dmm_tlbl_idx,
   input [CONFIG_DW-1:0]               msr_dmm_tlbl_nxt,
   input                               msr_dmm_tlbl_we,
   input [CONFIG_DTLB_P_SETS-1:0]      msr_dmm_tlbh_idx,
   input [CONFIG_DW-1:0]               msr_dmm_tlbh_nxt,
   input                               msr_dmm_tlbh_we
);
   localparam VPN_SHIFT                = CONFIG_P_PAGE_SIZE;
   localparam PPN_SHIFT                = VPN_SHIFT;
   localparam VPN_DW                   = CONFIG_AW-VPN_SHIFT;
   localparam PPN_DW                   = CONFIG_AW-PPN_SHIFT;
   assign msr_dmmid = {{32-3{1'b0}}, CONFIG_DTLB_P_SETS[2:0]};
   wire                                msr_psr_dmme_ff;
   wire                                msr_psr_rm_ff;
   wire                                we_ff;
   wire [VPN_DW-1:0]                   tgt_vpn_ff;
   wire [CONFIG_DW-1:0]                tlb_l_ff;
   wire [CONFIG_DW-1:0]                tlb_h_ff;
   wire [CONFIG_DTLB_P_SETS-1:0] tgt_index_nxt = vpn[CONFIG_DTLB_P_SETS-1:0];
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_dmme (.CLK(clk),.RST(rst), .LOAD(re), .D(msr_psr_dmme), .Q(msr_psr_dmme_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_rm (.CLK(clk),.RST(rst), .LOAD(re), .D(msr_psr_rm), .Q(msr_psr_rm_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_we (.CLK(clk),.RST(rst), .LOAD(re), .D(we), .Q(we_ff) );
   ysyx_20210479_mDFF_l #(.DW(VPN_DW)) ff_tgt_vpn (.CLK(clk), .LOAD(re), .D(vpn), .Q(tgt_vpn_ff) );
   ysyx_20210479_mRF_nwnr
      #(
         .DW      (CONFIG_DW),
         .AW      (CONFIG_DTLB_P_SETS),
         .NUM_READ (1),
         .NUM_WRITE (1)
      )
   U_TLB_L
      (
         .CLK     (clk),
         .RE      (re),
         .RADDR   (tgt_index_nxt),
         .RDATA   (tlb_l_ff),
         .WE      (msr_dmm_tlbl_we),
         .WADDR   (msr_dmm_tlbl_idx),
         .WDATA   (msr_dmm_tlbl_nxt)
      );
   ysyx_20210479_mRF_nwnr
      #(
         .DW      (CONFIG_DW),
         .AW      (CONFIG_DTLB_P_SETS),
         .NUM_READ (1),
         .NUM_WRITE (1)
      )
   U_TLB_H
      (
         .CLK     (clk),
         .RE      (re),
         .RADDR   (tgt_index_nxt),
         .RDATA   (tlb_h_ff),
         .WE      (msr_dmm_tlbh_we),
         .WADDR   (msr_dmm_tlbh_idx),
         .WDATA   (msr_dmm_tlbh_nxt)
      );
   wire tlb_v = tlb_l_ff[0];
   wire [VPN_DW-1:0] tlb_vpn = tlb_l_ff[CONFIG_DW-1:CONFIG_DW-VPN_DW];
   wire tlb_p = tlb_h_ff[0];
   wire tlb_uw = tlb_h_ff[3];
   wire tlb_ur = tlb_h_ff[4];
   wire tlb_rw = tlb_h_ff[5];
   wire tlb_rr = tlb_h_ff[6];
   wire tlb_unc = tlb_h_ff[7];
   wire tlb_s = tlb_h_ff[8];
   wire [PPN_DW-1:0] tlb_ppn = tlb_h_ff[CONFIG_DW-1:CONFIG_DW-PPN_DW];
   wire perm_denied;
   wire tlb_miss;
   assign perm_denied =
      (
         (msr_psr_rm_ff & ((we_ff & ~tlb_rw) | (~we_ff & ~tlb_rr)) ) |
         (~msr_psr_rm_ff & ((we_ff & ~tlb_uw) | (~we_ff & ~tlb_ur)) )
       );
   assign tlb_miss = ~(tlb_v & (tlb_vpn == tgt_vpn_ff));
   assign EDTM = tlb_miss & msr_psr_dmme_ff;
   assign EDPF = perm_denied & ~tlb_miss & msr_psr_dmme_ff;
   assign ppn = msr_psr_dmme_ff ? tlb_ppn : tgt_vpn_ff;
generate
   if (CONFIG_DMMU_ENABLE_UNCACHED_SEG)
      assign uncached = (msr_psr_dmme_ff & ~tlb_miss & ~perm_denied & tlb_unc) | (~EDTM & ~EDPF & ~ppn[CONFIG_AW-CONFIG_P_PAGE_SIZE-1]);
   else
      assign uncached = (msr_psr_dmme_ff & ~tlb_miss & ~perm_denied & tlb_unc);
endgenerate
endmodule
module ysyx_20210479_ex
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_DW = 0,
   parameter                           CONFIG_P_ISSUE_WIDTH = 0,
   parameter                           CONFIG_PHT_P_NUM = 0,
   parameter                           CONFIG_BTB_P_NUM = 0,
   parameter                           CONFIG_ENABLE_MUL = 0,
   parameter                           CONFIG_ENABLE_DIV = 0,
   parameter                           CONFIG_ENABLE_DIVU = 0,
   parameter                           CONFIG_ENABLE_MOD = 0,
   parameter                           CONFIG_ENABLE_MODU = 0,
   parameter                           CONFIG_ENABLE_ASR = 0,
   parameter                           CONFIG_NUM_IRQ = 0,
   parameter                           CONFIG_DC_P_WAYS = 0,
   parameter                           CONFIG_DC_P_SETS = 0,
   parameter                           CONFIG_DC_P_LINE = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_DMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_ITLB_P_SETS = 0,
   parameter                           CONFIG_DTLB_P_SETS = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EITM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_ESYSCALL_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EINSN_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIRQ_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDTM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EALIGN_VECTOR = 0,
   parameter                           AXI_P_DW_BYTES    = 0,
   parameter                           AXI_ADDR_WIDTH    = 0,
   parameter                           AXI_ID_WIDTH      = 0,
   parameter                           AXI_USER_WIDTH    = 0
)
(
   input                               clk,
   input                               rst,
   output                              stall,
   output                              flush,
   output [(CONFIG_AW-2 )-1:0]                  flush_tgt,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_valid,
   input [9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_alu_opc_bus,
   input [5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lpu_opc_bus,
   input [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_epu_opc_bus,
   input [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bru_opc_bus,
   input [7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lsu_opc_bus,
   input [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bpu_upd,
   input [(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_pc,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_imm,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand1,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand2,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_waddr,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_we,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_dout,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_dout,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_dout,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_wdat,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_we,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_we,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_we,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_we,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_waddr,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_waddr,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_waddr,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_waddr,
   output                              ro_ex_s1_load0,
   output                              ro_ex_s2_load0,
   output                              ro_ex_s3_load0,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_wdat,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_waddr,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_we,
   output                              bpu_wb,
   output                              bpu_wb_is_bcc,
   output                              bpu_wb_is_breg,
   output                              bpu_wb_is_brel,
   output                              bpu_wb_taken,
   output [(CONFIG_AW-2 )-1:0]                  bpu_wb_pc,
   output [(CONFIG_AW-2 )-1:0]                  bpu_wb_npc_act,
   output [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]             bpu_wb_upd,
   input [CONFIG_NUM_IRQ-1:0]          irqs,
   output                              irq_async,
   output                              tsc_irq,
   output                              msr_psr_imme,
   output                              msr_psr_rm,
   output                              msr_psr_ice,
   input [CONFIG_DW-1:0]               msr_immid,
   output [CONFIG_ITLB_P_SETS-1:0]     msr_imm_tlbl_idx,
   output [CONFIG_DW-1:0]              msr_imm_tlbl_nxt,
   output                              msr_imm_tlbl_we,
   output [CONFIG_ITLB_P_SETS-1:0]     msr_imm_tlbh_idx,
   output [CONFIG_DW-1:0]              msr_imm_tlbh_nxt,
   output                              msr_imm_tlbh_we,
   input [CONFIG_DW-1:0]               msr_icid,
   output [CONFIG_DW-1:0]              msr_icinv_nxt,
   output                              msr_icinv_we,
   input                               msr_icinv_ready,
   input                               dbus_ARREADY,
   output                              dbus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_ARADDR,
   output [2:0]                        dbus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_ARID,
   output [AXI_USER_WIDTH-1:0]         dbus_ARUSER,
   output [7:0]                        dbus_ARLEN,
   output [2:0]                        dbus_ARSIZE,
   output [1:0]                        dbus_ARBURST,
   output                              dbus_ARLOCK,
   output [3:0]                        dbus_ARCACHE,
   output [3:0]                        dbus_ARQOS,
   output [3:0]                        dbus_ARREGION,
   output                              dbus_RREADY,
   input                               dbus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_RDATA,
   input  [1:0]                        dbus_RRESP,
   input                               dbus_RLAST,
   input  [AXI_ID_WIDTH-1:0]           dbus_RID,
   input  [AXI_USER_WIDTH-1:0]         dbus_RUSER,
   input                               dbus_AWREADY,
   output                              dbus_AWVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_AWADDR,
   output [2:0]                        dbus_AWPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_AWID,
   output [AXI_USER_WIDTH-1:0]         dbus_AWUSER,
   output [7:0]                        dbus_AWLEN,
   output [2:0]                        dbus_AWSIZE,
   output [1:0]                        dbus_AWBURST,
   output                              dbus_AWLOCK,
   output [3:0]                        dbus_AWCACHE,
   output [3:0]                        dbus_AWQOS,
   output [3:0]                        dbus_AWREGION,
   input                               dbus_WREADY,
   output                              dbus_WVALID,
   output [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_WDATA,
   output [(1<<AXI_P_DW_BYTES)-1:0]    dbus_WSTRB,
   output                              dbus_WLAST,
   output [AXI_USER_WIDTH-1:0]         dbus_WUSER,
   output                              dbus_BREADY,
   input                               dbus_BVALID,
   input [1:0]                         dbus_BRESP,
   input [AXI_ID_WIDTH-1:0]            dbus_BID,
   input [AXI_USER_WIDTH-1:0]          dbus_BUSER
);
   localparam IW                       = (1<<CONFIG_P_ISSUE_WIDTH);
   wire [CONFIG_DW-1:0] epu_dout;               
   wire                 epu_dout_valid;         
   wire                 epu_s2i_EALIGN;         
   wire                 epu_s2i_EDPF;           
   wire                 epu_s2i_EDTM;           
   wire [CONFIG_AW-1:0] epu_s2i_vaddr;          
   wire                 exc_flush;              
   wire [(CONFIG_AW-2 )-1:0]     exc_flush_tgt;          
   wire                 lsu_stall_req;          
   wire [CONFIG_DW-1:0] msr_coreid;             
   wire [CONFIG_DW-1:0] msr_cpuid;              
   wire [CONFIG_DW-1:0] msr_dcfls_nxt;          
   wire                 msr_dcfls_we;           
   wire [CONFIG_DW-1:0] msr_dcid;               
   wire [CONFIG_DW-1:0] msr_dcinv_nxt;          
   wire                 msr_dcinv_we;           
   wire [CONFIG_DTLB_P_SETS-1:0] msr_dmm_tlbh_idx;
   wire [CONFIG_DW-1:0] msr_dmm_tlbh_nxt;       
   wire                 msr_dmm_tlbh_we;        
   wire [CONFIG_DTLB_P_SETS-1:0] msr_dmm_tlbl_idx;
   wire [CONFIG_DW-1:0] msr_dmm_tlbl_nxt;       
   wire                 msr_dmm_tlbl_we;        
   wire [CONFIG_DW-1:0] msr_dmmid;              
   wire [CONFIG_DW-1:0] msr_elsa;               
   wire [CONFIG_DW-1:0] msr_elsa_nxt;           
   wire                 msr_elsa_we;            
   wire [CONFIG_DW-1:0] msr_epc;                
   wire [CONFIG_DW-1:0] msr_epc_nxt;            
   wire                 msr_epc_we;             
   wire [10-1:0] msr_epsr;            
   wire [10-1:0] msr_epsr_nxt;        
   wire                 msr_epsr_we;            
   wire [10-1:0] msr_psr;             
   wire                 msr_psr_dce;            
   wire                 msr_psr_dce_nxt;        
   wire                 msr_psr_dce_we;         
   wire                 msr_psr_dmme;           
   wire                 msr_psr_dmme_nxt;       
   wire                 msr_psr_dmme_we;        
   wire                 msr_psr_ice_nxt;        
   wire                 msr_psr_ice_we;         
   wire                 msr_psr_imme_nxt;       
   wire                 msr_psr_imme_we;        
   wire                 msr_psr_ire;            
   wire                 msr_psr_ire_nxt;        
   wire                 msr_psr_ire_we;         
   wire                 msr_psr_restore;        
   wire                 msr_psr_rm_nxt;         
   wire                 msr_psr_rm_we;          
   wire                 msr_psr_save;           
   wire [CONFIG_DW*4-1:0] msr_sr;    
   wire [CONFIG_DW-1:0] msr_sr_nxt;             
   wire [4-1:0] msr_sr_we;           
   wire [CONFIG_DW-1:0]                bru_dout;
   wire                                bru_dout_valid;
   wire                                p_ce_s1;
   wire                                p_ce_s2;
   wire                                p_ce_s3;
   wire                                ex_lsu_load0;
   wire                                add_s                         [IW-1:0];
   wire [CONFIG_DW-1:0]                add_sum                       [IW-1:0];
   wire                                add_carry                     [IW-1:0];
   wire                                add_overflow                  [IW-1:0];
   wire                                b_taken;
   wire [(CONFIG_AW-2 )-1:0]                    b_tgt;
   wire                                is_bcc, is_breg, is_brel;
   wire                                agu_en;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]               ex_bpu_upd_unpacked           [IW-1:0];
   wire [(CONFIG_AW-2 )-1:0]                    npc                           [IW-1:0];
   reg [IW-1:0]                        cmt_valid_msk;
   wire                                icinv_stall_req;
   wire                                p_ce_s1_no_icinv_stall;
   wire [IW-1:0]                       se_fail_vec;
   wire [(CONFIG_AW-2 )*IW-1:0]                 se_tgt_vec;
   wire                                se_fail;
   wire [(CONFIG_AW-2 )-1:0]                    se_tgt;
   wire                                se_flush;
   wire                                flush_s1;
   wire                                flush_s2;
   wire [IW-1:0]                       s1i_cmt_valid;
   wire [CONFIG_DW*IW-1:0]             s1i_rf_dout_1, s1i_rf_dout;
   wire [IW-1:0]                       s1i_rf_we;
   wire [CONFIG_DW*IW-1:0]             s1o_rf_dout;
   wire [5*IW-1:0]          s1o_rf_waddr;
   wire [IW-1:0]                       s1o_rf_we;
   wire                                s1o_lsu_load0;
   wire                                s1o_se_flush;
   wire [(CONFIG_AW-2 )-1:0]                    s1o_se_flush_tgt;
   wire [CONFIG_DW-1:0]                s2o_lsu_dout0;
   wire                                s2o_lsu_load0;
   wire [CONFIG_DW*IW-1:0]             s2o_rf_dout;
   wire [5*IW-1:0]          s2o_rf_waddr;
   wire [IW-1:0]                       s2o_rf_we;
   wire [CONFIG_DW*IW-1:0]             s3i_rf_wdat;
   genvar i;
   integer j;
   generate
      for(i=0;i<IW;i=i+1)
         begin : gen_alus
            assign ex_bpu_upd_unpacked[i] = ex_bpu_upd[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)];
            ysyx_20210479_ex_add
               #(
                 .CONFIG_DW             (CONFIG_DW))
            U_ADD
               (
                  .a                   (ex_operand1[i*CONFIG_DW +: CONFIG_DW]),
                  .b                   (((i==0) & agu_en) ? ex_imm[i*CONFIG_DW +: CONFIG_DW] : ex_operand2[i*CONFIG_DW +: CONFIG_DW]),
                  .s                   (add_s[i]),
                  .sum                 (add_sum[i]),
                  .carry               (add_carry[i]),
                  .overflow            (add_overflow[i])
               );
            ysyx_20210479_ex_alu
               #(
                 .CONFIG_DW             (CONFIG_DW),
                 .CONFIG_ENABLE_MUL     (CONFIG_ENABLE_MUL),
                 .CONFIG_ENABLE_DIV     (CONFIG_ENABLE_DIV),
                 .CONFIG_ENABLE_DIVU    (CONFIG_ENABLE_DIVU),
                 .CONFIG_ENABLE_MOD     (CONFIG_ENABLE_MOD),
                 .CONFIG_ENABLE_MODU    (CONFIG_ENABLE_MODU),
                 .CONFIG_ENABLE_ASR     (CONFIG_ENABLE_ASR))
            U_ALU
               (
                  .ex_alu_opc_bus      (ex_alu_opc_bus[i*9  +: 9 ]),
                  .ex_operand1         (ex_operand1[i*CONFIG_DW +: CONFIG_DW]),
                  .ex_operand2         (ex_operand2[i*CONFIG_DW +: CONFIG_DW]),
                  .add_sum             (add_sum[i]),
                  .alu_result          (s1i_rf_dout_1[i*CONFIG_DW +: CONFIG_DW])
               );
            if (i > 0) 
               begin
                  assign add_s[i] = ex_alu_opc_bus[i*9  + 1];
                  assign s1i_rf_dout[i*CONFIG_DW +: CONFIG_DW] = s1i_rf_dout_1[i*CONFIG_DW +: CONFIG_DW];
               end
         end
   endgenerate
   ysyx_20210479_ex_bru
      #(
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_AW                      (CONFIG_AW))
   U_BRU
      (
         .ex_valid         (ex_valid[0]),
         .ex_bru_opc_bus   (ex_bru_opc_bus[0*8 +: 8]),
         .ex_pc            (ex_pc[0*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )]),
         .ex_imm           (ex_imm[0*CONFIG_DW +: CONFIG_DW]),
         .ex_operand1      (ex_operand1[0*CONFIG_DW +: CONFIG_DW]),
         .ex_operand2      (ex_operand2[0*CONFIG_DW +: CONFIG_DW]),
         .ex_rf_we         (ex_rf_we[0]),
         .npc              (npc[0]),
         .add_sum          (add_sum[0]),
         .add_carry        (add_carry[0]),
         .add_overflow     (add_overflow[0]),
         .b_taken          (b_taken),
         .b_tgt            (b_tgt),
         .is_bcc           (is_bcc),
         .is_breg          (is_breg),
         .is_brel          (is_brel),
         .bru_dout         (bru_dout),
         .bru_dout_valid   (bru_dout_valid)
      );
   ysyx_20210479_ex_epu
      #(
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_EITM_VECTOR             (CONFIG_EITM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIPF_VECTOR             (CONFIG_EIPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_ESYSCALL_VECTOR         (CONFIG_ESYSCALL_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EINSN_VECTOR            (CONFIG_EINSN_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIRQ_VECTOR             (CONFIG_EIRQ_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDTM_VECTOR             (CONFIG_EDTM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDPF_VECTOR             (CONFIG_EDPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EALIGN_VECTOR           (CONFIG_EALIGN_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_ITLB_P_SETS             (CONFIG_ITLB_P_SETS),
        .CONFIG_DTLB_P_SETS             (CONFIG_DTLB_P_SETS),
        .CONFIG_NUM_IRQ                 (CONFIG_NUM_IRQ))
   U_EPU
      (
       .epu_dout                        (epu_dout[CONFIG_DW-1:0]),
       .epu_dout_valid                  (epu_dout_valid),
       .exc_flush                       (exc_flush),
       .exc_flush_tgt                   (exc_flush_tgt[(CONFIG_AW-2 )-1:0]),
       .irq_async                       (irq_async),
       .tsc_irq                         (tsc_irq),
       .msr_psr_rm_nxt                  (msr_psr_rm_nxt),
       .msr_psr_rm_we                   (msr_psr_rm_we),
       .msr_psr_imme_nxt                (msr_psr_imme_nxt),
       .msr_psr_imme_we                 (msr_psr_imme_we),
       .msr_psr_dmme_nxt                (msr_psr_dmme_nxt),
       .msr_psr_dmme_we                 (msr_psr_dmme_we),
       .msr_psr_ire_nxt                 (msr_psr_ire_nxt),
       .msr_psr_ire_we                  (msr_psr_ire_we),
       .msr_psr_ice_nxt                 (msr_psr_ice_nxt),
       .msr_psr_ice_we                  (msr_psr_ice_we),
       .msr_psr_dce_nxt                 (msr_psr_dce_nxt),
       .msr_psr_dce_we                  (msr_psr_dce_we),
       .msr_psr_save                    (msr_psr_save),
       .msr_psr_restore                 (msr_psr_restore),
       .msr_epc_nxt                     (msr_epc_nxt[CONFIG_DW-1:0]),
       .msr_epc_we                      (msr_epc_we),
       .msr_epsr_nxt                    (msr_epsr_nxt[10-1:0]),
       .msr_epsr_we                     (msr_epsr_we),
       .msr_elsa_nxt                    (msr_elsa_nxt[CONFIG_DW-1:0]),
       .msr_elsa_we                     (msr_elsa_we),
       .msr_imm_tlbl_idx                (msr_imm_tlbl_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbl_nxt                (msr_imm_tlbl_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbl_we                 (msr_imm_tlbl_we),
       .msr_imm_tlbh_idx                (msr_imm_tlbh_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbh_nxt                (msr_imm_tlbh_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbh_we                 (msr_imm_tlbh_we),
       .msr_dmm_tlbl_idx                (msr_dmm_tlbl_idx[CONFIG_DTLB_P_SETS-1:0]),
       .msr_dmm_tlbl_nxt                (msr_dmm_tlbl_nxt[CONFIG_DW-1:0]),
       .msr_dmm_tlbl_we                 (msr_dmm_tlbl_we),
       .msr_dmm_tlbh_idx                (msr_dmm_tlbh_idx[CONFIG_DTLB_P_SETS-1:0]),
       .msr_dmm_tlbh_nxt                (msr_dmm_tlbh_nxt[CONFIG_DW-1:0]),
       .msr_dmm_tlbh_we                 (msr_dmm_tlbh_we),
       .msr_icinv_nxt                   (msr_icinv_nxt[CONFIG_DW-1:0]),
       .msr_icinv_we                    (msr_icinv_we),
       .msr_dcinv_nxt                   (msr_dcinv_nxt[CONFIG_DW-1:0]),
       .msr_dcinv_we                    (msr_dcinv_we),
       .msr_dcfls_nxt                   (msr_dcfls_nxt[CONFIG_DW-1:0]),
       .msr_dcfls_we                    (msr_dcfls_we),
       .msr_sr_nxt                      (msr_sr_nxt[CONFIG_DW-1:0]),
       .msr_sr_we                       (msr_sr_we[4-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .flush_s1                        (flush_s1),
       .p_ce_s1                         (p_ce_s1),
       .p_ce_s1_no_icinv_stall          (p_ce_s1_no_icinv_stall),
       .p_ce_s2                         (p_ce_s2),
       .ex_pc                           (ex_pc[0*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )]), 
       .ex_npc                          (npc[0]),                
       .ex_valid                        (s1i_cmt_valid[0]),      
       .ex_epu_opc_bus                  (ex_epu_opc_bus[0*8 +: 8]), 
       .ex_operand1                     (ex_operand1[0*CONFIG_DW +: CONFIG_DW]), 
       .ex_operand2                     (ex_operand2[0*CONFIG_DW +: CONFIG_DW]), 
       .ex_imm                          (ex_imm[0*CONFIG_DW +: CONFIG_DW]), 
       .s2i_EDTM                        (epu_s2i_EDTM),          
       .s2i_EDPF                        (epu_s2i_EDPF),          
       .s2i_EALIGN                      (epu_s2i_EALIGN),        
       .s2i_vaddr                       (epu_s2i_vaddr[CONFIG_AW-1:0]), 
       .irqs                            (irqs[CONFIG_NUM_IRQ-1:0]),
       .msr_psr                         (msr_psr[10-1:0]),
       .msr_psr_ire                     (msr_psr_ire),
       .msr_cpuid                       (msr_cpuid[CONFIG_DW-1:0]),
       .msr_epc                         (msr_epc[CONFIG_DW-1:0]),
       .msr_epsr                        (msr_epsr[10-1:0]),
       .msr_elsa                        (msr_elsa[CONFIG_DW-1:0]),
       .msr_coreid                      (msr_coreid[CONFIG_DW-1:0]),
       .msr_immid                       (msr_immid[CONFIG_DW-1:0]),
       .msr_dmmid                       (msr_dmmid[CONFIG_DW-1:0]),
       .msr_icid                        (msr_icid[CONFIG_DW-1:0]),
       .msr_dcid                        (msr_dcid[CONFIG_DW-1:0]),
       .msr_sr                          (msr_sr[CONFIG_DW*4-1:0]));
   assign add_s[0] =
      (
         ex_alu_opc_bus[0*9  + 1] |
         ex_bru_opc_bus[0*8 + 0] |
         ex_bru_opc_bus[0*8 + 1] |
         ex_bru_opc_bus[0*8 + 3] |
         ex_bru_opc_bus[0*8 + 2] |
         ex_bru_opc_bus[0*8 + 5] |
         ex_bru_opc_bus[0*8 + 4]
      );
   assign s1i_rf_dout[0*CONFIG_DW +: CONFIG_DW] =
      (epu_dout_valid)
         ? epu_dout
         : (bru_dout_valid)
            ? bru_dout
            : s1i_rf_dout_1[0*CONFIG_DW +: CONFIG_DW];
   ysyx_20210479_ex_lsu
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_DW                    (CONFIG_P_DW),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_DMMU_ENABLE_UNCACHED_SEG(CONFIG_DMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_DTLB_P_SETS             (CONFIG_DTLB_P_SETS),
        .CONFIG_DC_P_LINE               (CONFIG_DC_P_LINE),
        .CONFIG_DC_P_SETS               (CONFIG_DC_P_SETS),
        .CONFIG_DC_P_WAYS               (CONFIG_DC_P_WAYS),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_LSU
      (
       .lsu_stall_req                   (lsu_stall_req),
       .agu_en                          (agu_en),
       .dbus_ARVALID                    (dbus_ARVALID),
       .dbus_ARADDR                     (dbus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_ARPROT                     (dbus_ARPROT[2:0]),
       .dbus_ARID                       (dbus_ARID[AXI_ID_WIDTH-1:0]),
       .dbus_ARUSER                     (dbus_ARUSER[AXI_USER_WIDTH-1:0]),
       .dbus_ARLEN                      (dbus_ARLEN[7:0]),
       .dbus_ARSIZE                     (dbus_ARSIZE[2:0]),
       .dbus_ARBURST                    (dbus_ARBURST[1:0]),
       .dbus_ARLOCK                     (dbus_ARLOCK),
       .dbus_ARCACHE                    (dbus_ARCACHE[3:0]),
       .dbus_ARQOS                      (dbus_ARQOS[3:0]),
       .dbus_ARREGION                   (dbus_ARREGION[3:0]),
       .dbus_RREADY                     (dbus_RREADY),
       .dbus_AWVALID                    (dbus_AWVALID),
       .dbus_AWADDR                     (dbus_AWADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_AWPROT                     (dbus_AWPROT[2:0]),
       .dbus_AWID                       (dbus_AWID[AXI_ID_WIDTH-1:0]),
       .dbus_AWUSER                     (dbus_AWUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWLEN                      (dbus_AWLEN[7:0]),
       .dbus_AWSIZE                     (dbus_AWSIZE[2:0]),
       .dbus_AWBURST                    (dbus_AWBURST[1:0]),
       .dbus_AWLOCK                     (dbus_AWLOCK),
       .dbus_AWCACHE                    (dbus_AWCACHE[3:0]),
       .dbus_AWQOS                      (dbus_AWQOS[3:0]),
       .dbus_AWREGION                   (dbus_AWREGION[3:0]),
       .dbus_WVALID                     (dbus_WVALID),
       .dbus_WDATA                      (dbus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_WSTRB                      (dbus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]),
       .dbus_WLAST                      (dbus_WLAST),
       .dbus_WUSER                      (dbus_WUSER[AXI_USER_WIDTH-1:0]),
       .dbus_BREADY                     (dbus_BREADY),
       .lsu_EDTM                        (epu_s2i_EDTM),          
       .lsu_EDPF                        (epu_s2i_EDPF),          
       .lsu_EALIGN                      (epu_s2i_EALIGN),        
       .lsu_vaddr                       (epu_s2i_vaddr[CONFIG_AW-1:0]), 
       .lsu_dout                        (s2o_lsu_dout0),         
       .msr_dmmid                       (msr_dmmid[CONFIG_DW-1:0]),
       .msr_dcid                        (msr_dcid[CONFIG_DW-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .p_ce_s1                         (p_ce_s1),
       .flush_s1                        (flush_s1),
       .ex_valid                        (s1i_cmt_valid[0]),      
       .ex_lsu_opc_bus                  (ex_lsu_opc_bus[0*7 +: 7]), 
       .add_sum                         (add_sum[0]),            
       .ex_operand2                     (ex_operand2[0*CONFIG_DW +: CONFIG_DW]), 
       .dbus_ARREADY                    (dbus_ARREADY),
       .dbus_RVALID                     (dbus_RVALID),
       .dbus_RDATA                      (dbus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_RRESP                      (dbus_RRESP[1:0]),
       .dbus_RLAST                      (dbus_RLAST),
       .dbus_RID                        (dbus_RID[AXI_ID_WIDTH-1:0]),
       .dbus_RUSER                      (dbus_RUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWREADY                    (dbus_AWREADY),
       .dbus_WREADY                     (dbus_WREADY),
       .dbus_BVALID                     (dbus_BVALID),
       .dbus_BRESP                      (dbus_BRESP[1:0]),
       .dbus_BID                        (dbus_BID[AXI_ID_WIDTH-1:0]),
       .dbus_BUSER                      (dbus_BUSER[AXI_USER_WIDTH-1:0]),
       .msr_psr_dmme                    (msr_psr_dmme),
       .msr_psr_rm                      (msr_psr_rm),
       .msr_psr_dce                     (msr_psr_dce),
       .msr_dmm_tlbl_idx                (msr_dmm_tlbl_idx[CONFIG_DTLB_P_SETS-1:0]),
       .msr_dmm_tlbl_nxt                (msr_dmm_tlbl_nxt[CONFIG_DW-1:0]),
       .msr_dmm_tlbl_we                 (msr_dmm_tlbl_we),
       .msr_dmm_tlbh_idx                (msr_dmm_tlbh_idx[CONFIG_DTLB_P_SETS-1:0]),
       .msr_dmm_tlbh_nxt                (msr_dmm_tlbh_nxt[CONFIG_DW-1:0]),
       .msr_dmm_tlbh_we                 (msr_dmm_tlbh_we),
       .msr_dcinv_nxt                   (msr_dcinv_nxt[CONFIG_DW-1:0]),
       .msr_dcinv_we                    (msr_dcinv_we),
       .msr_dcfls_nxt                   (msr_dcfls_nxt[CONFIG_DW-1:0]),
       .msr_dcfls_we                    (msr_dcfls_we));
   ysyx_20210479_ex_psr
      #(
        .CONFIG_DW                      (CONFIG_DW),
        .CPUID_VER                      (1),
        .CPUID_REV                      (0),
        .CPUID_FIMM                     (1),
        .CPUID_FDMM                     (1),
        .CPUID_FICA                     (1),
        .CPUID_FDCA                     (1),
        .CPUID_FDBG                     (0),
        .CPUID_FFPU                     (0),
        .CPUID_FIRQC                    (1),
        .CPUID_FTSC                     (1)
     )
   U_PSR
      (
       .msr_psr                         (msr_psr[10-1:0]),
       .msr_psr_rm                      (msr_psr_rm),
       .msr_psr_ire                     (msr_psr_ire),
       .msr_psr_imme                    (msr_psr_imme),
       .msr_psr_dmme                    (msr_psr_dmme),
       .msr_psr_ice                     (msr_psr_ice),
       .msr_psr_dce                     (msr_psr_dce),
       .msr_cpuid                       (msr_cpuid[CONFIG_DW-1:0]),
       .msr_epsr                        (msr_epsr[10-1:0]),
       .msr_epc                         (msr_epc[CONFIG_DW-1:0]),
       .msr_elsa                        (msr_elsa[CONFIG_DW-1:0]),
       .msr_coreid                      (msr_coreid[CONFIG_DW-1:0]),
       .msr_sr                          (msr_sr[CONFIG_DW*4-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .msr_psr_save                    (msr_psr_save),
       .msr_psr_restore                 (msr_psr_restore),
       .msr_psr_rm_nxt                  (msr_psr_rm_nxt),
       .msr_psr_rm_we                   (msr_psr_rm_we),
       .msr_psr_ire_nxt                 (msr_psr_ire_nxt),
       .msr_psr_ire_we                  (msr_psr_ire_we),
       .msr_psr_imme_nxt                (msr_psr_imme_nxt),
       .msr_psr_imme_we                 (msr_psr_imme_we),
       .msr_psr_dmme_nxt                (msr_psr_dmme_nxt),
       .msr_psr_dmme_we                 (msr_psr_dmme_we),
       .msr_psr_ice_nxt                 (msr_psr_ice_nxt),
       .msr_psr_ice_we                  (msr_psr_ice_we),
       .msr_psr_dce_nxt                 (msr_psr_dce_nxt),
       .msr_psr_dce_we                  (msr_psr_dce_we),
       .msr_epsr_nxt                    (msr_epsr_nxt[10-1:0]),
       .msr_epsr_we                     (msr_epsr_we),
       .msr_epc_nxt                     (msr_epc_nxt[CONFIG_DW-1:0]),
       .msr_epc_we                      (msr_epc_we),
       .msr_elsa_nxt                    (msr_elsa_nxt[CONFIG_DW-1:0]),
       .msr_elsa_we                     (msr_elsa_we),
       .msr_sr_nxt                      (msr_sr_nxt[CONFIG_DW-1:0]),
       .msr_sr_we                       (msr_sr_we[4-1:0]));
   generate
      for(i=0;i<IW;i=i+1)
         assign npc[i] = (ex_pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )]+'b1);
   endgenerate
   assign se_fail_vec[0] = ex_valid[0] & ((b_taken ^ ex_bpu_upd_unpacked[0][0]) | (b_tgt != ex_bpu_upd_unpacked[0][(CONFIG_AW-2 ):1])); 
   assign se_tgt_vec[0 +: (CONFIG_AW-2 )] = (b_taken) ? b_tgt : npc[0];
   generate
      for(i=1;i<IW;i=i+1)
         begin
            assign se_fail_vec[i] = ex_valid[i] & (1'b0 ^ ex_bpu_upd_unpacked[i][0]);
            assign se_tgt_vec[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )] = npc[i];
         end
   endgenerate
   ysyx_20210479_pmux_v #(.SELW(IW), .DW((CONFIG_AW-2 ))) pmux_se_tgt (.sel(se_fail_vec), .din(se_tgt_vec), .dout(se_tgt), .valid(se_fail) );
   always @(*)
      begin
         cmt_valid_msk[0] = 'b1;
         for(j=1;j<IW;j=j+1)
            cmt_valid_msk[j] = cmt_valid_msk[j-1] & ~se_fail_vec[j-1];
      end
   assign s1i_cmt_valid = (ex_valid & cmt_valid_msk);
   assign se_flush = (s1o_se_flush & p_ce_s2);
   assign bpu_wb = ex_valid[0];
   assign bpu_wb_is_bcc = is_bcc;
   assign bpu_wb_is_breg = is_breg;
   assign bpu_wb_is_brel = is_brel;
   assign bpu_wb_taken = b_taken;
   assign bpu_wb_pc = ex_pc[0 +: (CONFIG_AW-2 )];
   assign bpu_wb_npc_act = se_tgt_vec[0 +: (CONFIG_AW-2 )];
   assign bpu_wb_upd = ex_bpu_upd[0*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)];
   assign s1i_rf_we = (s1i_cmt_valid & ex_rf_we);
   assign s3i_rf_wdat[0 +: CONFIG_DW] = (s2o_lsu_load0)
                                          ? s2o_lsu_dout0
                                          : s2o_rf_dout[0 +: CONFIG_DW];
   generate
      for(i=1;i<IW;i=i+1)
         assign s3i_rf_wdat[i*CONFIG_DW +: CONFIG_DW] = s2o_rf_dout[i*CONFIG_DW +: CONFIG_DW];
   endgenerate
   assign ex_lsu_load0 = ex_lsu_opc_bus[0*7 + 0];
   assign ro_ex_s1_rf_dout = s1i_rf_dout;
   assign ro_ex_s2_rf_dout = s1o_rf_dout;
   assign ro_ex_s3_rf_dout = s2o_rf_dout;
   assign ro_cmt_rf_wdat = commit_rf_wdat;
   assign ro_ex_s1_rf_we = s1i_rf_we;
   assign ro_ex_s2_rf_we = s1o_rf_we;
   assign ro_ex_s3_rf_we = s2o_rf_we;
   assign ro_cmt_rf_we = commit_rf_we;
   assign ro_ex_s1_rf_waddr = ex_rf_waddr;
   assign ro_ex_s2_rf_waddr = s1o_rf_waddr;
   assign ro_ex_s3_rf_waddr = s2o_rf_waddr;
   assign ro_cmt_rf_waddr = commit_rf_waddr;
   assign ro_ex_s1_load0 = ex_lsu_load0;
   assign ro_ex_s2_load0 = s1o_lsu_load0;
   assign ro_ex_s3_load0 = s2o_lsu_load0;
   assign icinv_stall_req = (msr_icinv_we & ~msr_icinv_ready);
   assign stall = (lsu_stall_req | icinv_stall_req | 1'b0);
   assign p_ce_s1 = (p_ce_s1_no_icinv_stall & ~icinv_stall_req);
   assign p_ce_s1_no_icinv_stall = ~(lsu_stall_req | 1'b0);
   assign p_ce_s2 = ~(lsu_stall_req);
   assign p_ce_s3 = ~(lsu_stall_req);
   assign flush_s1 = (exc_flush | se_flush);
   assign flush_s2 = (exc_flush);
   assign flush = (exc_flush | se_flush);
   assign flush_tgt = (exc_flush)
                        ? exc_flush_tgt
                        : s1o_se_flush_tgt; 
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_se_flush (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(se_fail & ~flush_s1), .Q(s1o_se_flush) );
   ysyx_20210479_mDFF_l # (.DW((CONFIG_AW-2 ))) ff_s1o_se_flush_tgt (.CLK(clk), .LOAD(p_ce_s1), .D(se_tgt), .Q(s1o_se_flush_tgt) );
   ysyx_20210479_mDFF_l # (.DW(5*IW)) ff_s1o_rf_waddr (.CLK(clk), .LOAD(p_ce_s1), .D(ex_rf_waddr), .Q(s1o_rf_waddr) );
   ysyx_20210479_mDFF_lr # (.DW(IW)) ff_s1o_rf_we (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_rf_we & {IW{~flush_s1}}), .Q(s1o_rf_we) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW*IW)) ff_s1o_rf_dout (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_rf_dout), .Q(s1o_rf_dout) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_lsu_load (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(ex_lsu_load0 & ~flush_s1), .Q(s1o_lsu_load0) );
   ysyx_20210479_mDFF_l # (.DW(5*IW)) ff_s2o_rf_waddr (.CLK(clk), .LOAD(p_ce_s2), .D(s1o_rf_waddr), .Q(s2o_rf_waddr) );
   ysyx_20210479_mDFF_lr # (.DW(IW)) ff_s2o_rf_we (.CLK(clk), .RST(rst), .LOAD(p_ce_s2|flush_s2), .D(s1o_rf_we & {IW{~flush_s2}}), .Q(s2o_rf_we) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW*IW)) ff_s2o_rf_dout (.CLK(clk), .LOAD(p_ce_s2), .D(s1o_rf_dout), .Q(s2o_rf_dout) );
   ysyx_20210479_mDFF_l # (.DW(1)) ff_s2o_lsu_load (.CLK(clk), .LOAD(p_ce_s2), .D(s1o_lsu_load0), .Q(s2o_lsu_load0) );
   ysyx_20210479_mDFF_l # (.DW(5*IW)) ff_commit_rf_waddr (.CLK(clk), .LOAD(p_ce_s3), .D(s2o_rf_waddr), .Q(commit_rf_waddr) );
   ysyx_20210479_mDFF_lr # (.DW(IW)) ff_commit_rf_we (.CLK(clk), .RST(rst), .LOAD(p_ce_s3), .D(s2o_rf_we), .Q(commit_rf_we) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW*IW)) ff_commit_rf_wdat (.CLK(clk), .LOAD(p_ce_s3), .D(s3i_rf_wdat), .Q(commit_rf_wdat) );
endmodule
module ysyx_20210479_ex_add
#(
   parameter                           CONFIG_DW = 0
)
(
   input [CONFIG_DW-1:0]               a,
   input [CONFIG_DW-1:0]               b,
   input                               s,
   output [CONFIG_DW-1:0]              sum,
   output                              carry,
   output                              overflow
);
   wire                                ci;
   wire [CONFIG_DW-1:0]                op2;
   assign op2 = (s) ? ~b : b;
   assign ci = (s);
   assign {carry, sum} = a + op2 + {{CONFIG_DW-1{1'b0}}, ci};
   assign overflow = ((a[CONFIG_DW-1] == op2[CONFIG_DW-1]) &
                        (a[CONFIG_DW-1] ^ sum[CONFIG_DW-1]));
endmodule
module ysyx_20210479_ex_alu
#(
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_ENABLE_MUL = 0,
   parameter                           CONFIG_ENABLE_DIV = 0,
   parameter                           CONFIG_ENABLE_DIVU = 0,
   parameter                           CONFIG_ENABLE_MOD = 0,
   parameter                           CONFIG_ENABLE_MODU = 0,
   parameter                           CONFIG_ENABLE_ASR = 0
)
(
   input [9 -1:0]          ex_alu_opc_bus,
   input [CONFIG_DW-1:0]               ex_operand1,
   input [CONFIG_DW-1:0]               ex_operand2,
   input [CONFIG_DW-1:0]               add_sum,
   output [CONFIG_DW-1:0]              alu_result
);
   wire [CONFIG_DW-1:0]                dat_adder;
   wire [CONFIG_DW-1:0]                dat_and;
   wire [CONFIG_DW-1:0]                dat_or;
   wire [CONFIG_DW-1:0]                dat_xor;
   wire [CONFIG_DW-1:0]                dat_shifter;
   wire [CONFIG_DW-1:0]                dat_move;
   wire                                sel_adder;
   wire                                sel_and;
   wire                                sel_or;
   wire                                sel_xor;
   wire                                sel_shifter;
   wire                                sel_move;
   assign dat_adder = add_sum;
   assign sel_adder = (ex_alu_opc_bus[0] | ex_alu_opc_bus[1]);
   assign dat_and = (ex_operand1 & ex_operand2);
   assign dat_or = (ex_operand1 | ex_operand2);
   assign dat_xor = (ex_operand1 ^ ex_operand2);
   assign sel_and = ex_alu_opc_bus[3];
   assign sel_or = ex_alu_opc_bus[4];
   assign sel_xor = ex_alu_opc_bus[5];
   wire [CONFIG_DW-1:0] shift_right;
   wire [CONFIG_DW-1:0] shift_lsw;
   function [CONFIG_DW-1:0] reverse_bits;
      input [CONFIG_DW-1:0] a;
	   integer 			       i;
	   begin
         for(i=0; i<CONFIG_DW; i=i+1)
            reverse_bits[CONFIG_DW-1-i] = a[i];
      end
   endfunction
   assign shift_lsw = ex_alu_opc_bus[6] ? reverse_bits(ex_operand1) : ex_operand1;
   generate
      if (CONFIG_ENABLE_ASR)
         begin : gen_asr
            wire [CONFIG_DW-1:0] shift_msw;
            wire [CONFIG_DW*2-1:0] shift_wide;
            assign shift_msw = ex_alu_opc_bus[8] ? {CONFIG_DW{ex_operand1[CONFIG_DW-1]}} : {CONFIG_DW{1'b0}};
            assign shift_wide = {shift_msw, shift_lsw} >> ex_operand2[4:0];
            assign shift_right = shift_wide[CONFIG_DW-1:0];
         end
      else
         assign shift_right = shift_lsw >> ex_operand2[4:0];
   endgenerate
   assign dat_shifter = ex_alu_opc_bus[6] ? reverse_bits(shift_right) : shift_right;
   assign sel_shifter = ex_alu_opc_bus[6] | ex_alu_opc_bus[7] | ex_alu_opc_bus[8];
   assign sel_move = ex_alu_opc_bus[2];
   assign dat_move = {ex_operand2[16:0], 15'b0};
   assign alu_result =
      ({CONFIG_DW{sel_adder}} & dat_adder) |
      ({CONFIG_DW{sel_and}} & dat_and) |
      ({CONFIG_DW{sel_or}} & dat_or) |
      ({CONFIG_DW{sel_xor}} & dat_xor) |
      ({CONFIG_DW{sel_shifter}} & dat_shifter) |
      ({CONFIG_DW{sel_move}} & dat_move);
endmodule
module ysyx_20210479_ex_bru
#(
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_AW = 0
)
(
   input                               ex_valid,
   input [8-1:0]          ex_bru_opc_bus,
   input [(CONFIG_AW-2 )-1:0]                   ex_pc,
   input [CONFIG_DW-1:0]               ex_imm,
   input [CONFIG_DW-1:0]               ex_operand1,
   input [CONFIG_DW-1:0]               ex_operand2,
   input                               ex_rf_we,
   input [(CONFIG_AW-2 )-1:0]                   npc,
   input [CONFIG_DW-1:0]               add_sum,
   input                               add_carry,
   input                               add_overflow,
   output                              b_taken,
   output [(CONFIG_AW-2 )-1:0]                  b_tgt,
   output                              is_bcc,
   output                              is_breg,
   output                              is_brel,
   output [CONFIG_DW-1:0]              bru_dout,
   output                              bru_dout_valid
);
   wire                                cmp_eq;
   wire                                cmp_lt_s;
   wire                                cmp_lt_u;
   wire                                bcc_taken;
   wire                                b_lnk;
   assign cmp_eq = (ex_operand1 == ex_operand2);
   assign cmp_lt_s = (add_sum[CONFIG_DW-1] ^ add_overflow);
   assign cmp_lt_u = ~add_carry;
   assign is_bcc = (ex_bru_opc_bus[0] |
                     ex_bru_opc_bus[1] |
                     ex_bru_opc_bus[3] |
                     ex_bru_opc_bus[2] |
                     ex_bru_opc_bus[5] |
                     ex_bru_opc_bus[4]);
   assign is_breg = (ex_bru_opc_bus[6]);
   assign is_brel = (ex_bru_opc_bus[7]);
   assign bcc_taken = (ex_bru_opc_bus[0] & cmp_eq) |
                        (ex_bru_opc_bus[1] & ~cmp_eq) |
                        (ex_bru_opc_bus[3] & (~cmp_lt_u & ~cmp_eq)) |
                        (ex_bru_opc_bus[2] & (~cmp_lt_s & ~cmp_eq)) |
                        (ex_bru_opc_bus[5] & (cmp_lt_u | cmp_eq)) |
                        (ex_bru_opc_bus[4] & (cmp_lt_s | cmp_eq));
   assign b_taken = (ex_valid & (bcc_taken | is_breg | is_brel));
   assign b_tgt =
      ({(CONFIG_AW-2 ){bcc_taken}} & (ex_pc + ex_imm[CONFIG_AW-1:2 ])) |
      ({(CONFIG_AW-2 ){is_brel}} & (ex_pc + ex_operand2[CONFIG_AW-1:2 ])) |
      ({(CONFIG_AW-2 ){is_breg}} & ex_operand1[CONFIG_AW-1:2 ]);
   assign b_lnk = ((is_brel | is_breg) & ex_rf_we);
   assign bru_dout = {npc, {2 {1'b0}}};
   assign bru_dout_valid = b_lnk;
endmodule
module ysyx_20210479_ex_epu
#(
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_AW = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EITM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_ESYSCALL_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EINSN_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIRQ_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDTM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EALIGN_VECTOR = 0,
   parameter                           CONFIG_ITLB_P_SETS = 0,
   parameter                           CONFIG_DTLB_P_SETS = 0,
   parameter                           CONFIG_NUM_IRQ = 0
)
(
   input                               clk,
   input                               rst,
   input                               flush_s1,
   input                               p_ce_s1,
   input                               p_ce_s1_no_icinv_stall,
   input                               p_ce_s2,
   input [(CONFIG_AW-2 )-1:0]                   ex_pc,
   input [(CONFIG_AW-2 )-1:0]                   ex_npc,
   input                               ex_valid,
   input [8-1:0]          ex_epu_opc_bus,
   input [CONFIG_DW-1:0]               ex_operand1,
   input [CONFIG_DW-1:0]               ex_operand2,
   input [CONFIG_DW-1:0]               ex_imm,
   input                               s2i_EDTM,
   input                               s2i_EDPF,
   input                               s2i_EALIGN,
   input [CONFIG_AW-1:0]               s2i_vaddr,
   output [CONFIG_DW-1:0]              epu_dout,
   output                              epu_dout_valid,
   output                              exc_flush,
   output [(CONFIG_AW-2 )-1:0]                  exc_flush_tgt,
   input [CONFIG_NUM_IRQ-1:0]          irqs,
   output                              irq_async,
   output                              tsc_irq,
   input [10-1:0]            msr_psr,
   input                               msr_psr_ire,
   output                              msr_psr_rm_nxt,
   output                              msr_psr_rm_we,
   output                              msr_psr_imme_nxt,
   output                              msr_psr_imme_we,
   output                              msr_psr_dmme_nxt,
   output                              msr_psr_dmme_we,
   output                              msr_psr_ire_nxt,
   output                              msr_psr_ire_we,
   output                              msr_psr_ice_nxt,
   output                              msr_psr_ice_we,
   output                              msr_psr_dce_nxt,
   output                              msr_psr_dce_we,
   output                              msr_psr_save,
   output                              msr_psr_restore,
   input [CONFIG_DW-1:0]               msr_cpuid,
   input [CONFIG_DW-1:0]               msr_epc,
   output [CONFIG_DW-1:0]              msr_epc_nxt,
   output                              msr_epc_we,
   input [10-1:0]            msr_epsr,
   output [10-1:0]           msr_epsr_nxt,
   output                              msr_epsr_we,
   input [CONFIG_DW-1:0]               msr_elsa,
   output [CONFIG_DW-1:0]              msr_elsa_nxt,
   output                              msr_elsa_we,
   input [CONFIG_DW-1:0]               msr_coreid,
   input [CONFIG_DW-1:0]               msr_immid,
   output [CONFIG_ITLB_P_SETS-1:0]     msr_imm_tlbl_idx,
   output [CONFIG_DW-1:0]              msr_imm_tlbl_nxt,
   output                              msr_imm_tlbl_we,
   output [CONFIG_ITLB_P_SETS-1:0]     msr_imm_tlbh_idx,
   output [CONFIG_DW-1:0]              msr_imm_tlbh_nxt,
   output                              msr_imm_tlbh_we,
   input [CONFIG_DW-1:0]               msr_dmmid,
   output [CONFIG_DTLB_P_SETS-1:0]     msr_dmm_tlbl_idx,
   output [CONFIG_DW-1:0]              msr_dmm_tlbl_nxt,
   output                              msr_dmm_tlbl_we,
   output [CONFIG_DTLB_P_SETS-1:0]     msr_dmm_tlbh_idx,
   output [CONFIG_DW-1:0]              msr_dmm_tlbh_nxt,
   output                              msr_dmm_tlbh_we,
   input [CONFIG_DW-1:0]               msr_icid,
   output [CONFIG_DW-1:0]              msr_icinv_nxt,
   output                              msr_icinv_we,
   input [CONFIG_DW-1:0]               msr_dcid,
   output [CONFIG_DW-1:0]              msr_dcinv_nxt,
   output                              msr_dcinv_we,
   output [CONFIG_DW-1:0]              msr_dcfls_nxt,
   output                              msr_dcfls_we,
   input [CONFIG_DW*4-1:0]  msr_sr,
   output [CONFIG_DW-1:0]              msr_sr_nxt,
   output [4-1:0]           msr_sr_we
);
   localparam NCPU_WMSR_WE_W           = (12 + 9);
   wire [CONFIG_DW-1:0] msr_irqc_imr;           
   wire [CONFIG_DW-1:0] msr_irqc_irr;           
   wire [CONFIG_DW-1:0] msr_tsc_tcr;            
   wire [CONFIG_DW-1:0] msr_tsc_tsr;            
   wire [CONFIG_DW-1:0]                msr_irqc_imr_nxt;
   wire                                msr_irqc_imr_we;
   wire [CONFIG_DW-1:0]                msr_tsc_tsr_nxt;
   wire                                msr_tsc_tsr_we;
   wire [CONFIG_DW-1:0]                msr_tsc_tcr_nxt;
   wire                                msr_tsc_tcr_we;
   wire [CONFIG_DW-1:0]                s1i_msr_addr;
   wire [(14-9) -1:0]        s1i_bank_addr;
   wire [9-1:0]    s1i_bank_off;
   wire                                s1i_bank_ps;
   wire                                s1i_bank_imm;
   wire                                s1i_bank_dmm;
   wire                                s1i_bank_ic;
   wire                                s1i_bank_dc;
   wire                                s1i_bank_dbg;
   wire                                s1i_bank_irqc;
   wire                                s1i_bank_tsc;
   wire                                s1i_bank_sr;
   wire [CONFIG_DW-1:0]                dout_ps;
   wire                                msr_imm_tlbl_sel;
   wire                                msr_imm_tlbh_sel;
   wire [CONFIG_DW-1:0]                dout_imm;
   wire                                msr_dmm_tlbl_sel;
   wire                                msr_dmm_tlbh_sel;
   wire                                msr_ic_id_sel;
   wire                                msr_ic_inv_sel;
   wire                                msr_dc_id_sel;
   wire                                msr_dc_inv_sel;
   wire                                msr_dc_fls_sel;
   wire [CONFIG_DW-1:0]                dout_dmm;
   wire [CONFIG_DW-1:0]                dout_ic;
   wire [CONFIG_DW-1:0]                dout_dc;
   wire                                msr_irqc_imr_sel;
   wire                                msr_irqc_irr_sel;
   wire [CONFIG_DW-1:0]                dout_irqc;
   wire                                msr_tsc_tsr_sel;
   wire                                msr_tsc_tcr_sel;
   wire [CONFIG_DW-1:0]                dout_tsc;
   wire [CONFIG_DW-1:0]                dout_sr;
   wire                                s1i_wmsr_psr_we;
   wire                                s1i_wmsr_epc_we;
   wire                                s1i_wmsr_epsr_we;
   wire                                s1i_wmsr_elsa_we;
   wire                                s1i_msr_imm_tlbl_we;
   wire                                s1i_msr_imm_tlbh_we;
   wire                                s1i_msr_dmm_tlbl_we;
   wire                                s1i_msr_dmm_tlbh_we;
   wire                                s1i_msr_ic_inv_we;
   wire                                s1i_msr_dc_inv_we;
   wire                                s1i_msr_dc_fls_we;
   wire                                s1i_msr_irqc_imr_we;
   wire                                s1i_msr_tsc_tsr_we;
   wire                                s1i_msr_tsc_tcr_we;
   wire                                s1i_msr_sr_we;
   wire   [CONFIG_DW-1:0]              s1i_msr_wdat;
   wire   [NCPU_WMSR_WE_W-1:0]         s1i_wmsr_we;
   wire                                s1i_ERET;
   wire                                s1i_ESYSCALL;
   wire                                s1i_EINSN;
   wire                                s1i_EIPF;
   wire                                s1i_EITM;
   wire                                s1i_EIRQ;
   wire                                s1i_E_FLUSH_TLB;
   wire                                s1o_commit_wmsr_psr_we;
   wire                                s1o_commit_wmsr_epc_we;
   wire                                s1o_commit_wmsr_epsr_we;
   wire                                s1o_commit_wmsr_elsa_we;
   wire                                s1o_commit_msr_imm_tlbl_we;
   wire                                s1o_commit_msr_imm_tlbh_we;
   wire                                s1o_commit_msr_dmm_tlbl_we;
   wire                                s1o_commit_msr_dmm_tlbh_we;
   wire                                s1o_commit_msr_irqc_imr_we;
   wire                                s1o_commit_msr_tsc_tsr_we;
   wire                                s1o_commit_msr_tsc_tcr_we;
   wire                                s1o_commit_msr_sr_we;
   wire [9-1:0]    s1o_commit_bank_off;
   wire  [(CONFIG_AW-2 )-1:0]                   s1o_commit_epc;
   wire [(CONFIG_AW-2 )-1:0]                    s1o_commit_nepc;
   wire                                s1o_commit_ERET;
   wire                                s1o_commit_ESYSCALL;
   wire                                s1o_commit_EINSN;
   wire                                s1o_commit_EIPF;
   wire                                s1o_commit_EITM;
   wire                                s1o_commit_EIRQ;
   wire                                s1o_commit_E_FLUSH_TLB;
   wire  [NCPU_WMSR_WE_W-1:0]          s1o_commit_wmsr_we;
   wire  [CONFIG_DW-1:0]               s1o_commit_wmsr_dat;
   wire                                s1o_wmsr_psr_rm;
   wire                                s1o_wmsr_psr_ire;
   wire                                s1o_wmsr_psr_imme;
   wire                                s1o_wmsr_psr_dmme;
   wire                                s1o_wmsr_psr_ice;
   wire                                s1o_wmsr_psr_dce;
   wire                                s1o_set_elsa_as_pc;
   wire                                s1o_set_elsa;
   wire [CONFIG_DW-1:0]                s1o_lsa_nxt;
   genvar i;
   assign s1i_msr_wdat = ex_operand2;
   assign s1i_msr_addr = ex_operand1 | {{CONFIG_DW-15{1'b0}}, ex_imm[14:0]};
   assign s1i_bank_addr = s1i_msr_addr[(14-9) +9-1:9];
   assign s1i_bank_off = s1i_msr_addr[9-1:0];
   assign dout_ps =
      (
         ({CONFIG_DW{s1i_bank_off[0]}} & {{CONFIG_DW-10{1'b0}}, msr_psr[10-1:0]}) |
         ({CONFIG_DW{s1i_bank_off[1]}} & msr_cpuid) |
         ({CONFIG_DW{s1i_bank_off[2]}} & {{CONFIG_DW-10{1'b0}}, msr_epsr[10-1:0]}) |
         ({CONFIG_DW{s1i_bank_off[3]}} & msr_epc) |
         ({CONFIG_DW{s1i_bank_off[4]}} & msr_elsa) |
         ({CONFIG_DW{s1i_bank_off[5]}} & msr_coreid)
      );
   assign msr_imm_tlbl_sel = s1i_bank_off[8] & ~s1i_bank_off[7];
   assign msr_imm_tlbh_sel = s1i_bank_off[8] & s1i_bank_off[7];
   assign dout_imm =
      (
         ({CONFIG_DW{~s1i_bank_off[8]}} & msr_immid)
      );
   assign msr_dmm_tlbl_sel = s1i_bank_off[8] & ~s1i_bank_off[7];
   assign msr_dmm_tlbh_sel = s1i_bank_off[8] & s1i_bank_off[7];
   assign dout_dmm =
      (
         ({CONFIG_DW{~s1i_bank_off[8]}} & msr_dmmid)
      );
   assign msr_ic_id_sel = s1i_bank_off[0];
   assign msr_ic_inv_sel = s1i_bank_off[1];
   assign dout_ic =
      (
         ({CONFIG_DW{msr_ic_id_sel}} & msr_icid)
      );
   assign msr_dc_id_sel = s1i_bank_off[0];
   assign msr_dc_inv_sel = s1i_bank_off[1];
   assign msr_dc_fls_sel = s1i_bank_off[2];
   assign dout_dc =
      (
         ({CONFIG_DW{msr_dc_id_sel}} & msr_dcid)
      );
   assign msr_irqc_imr_sel = s1i_bank_off[0];
   assign msr_irqc_irr_sel = s1i_bank_off[1];
   assign dout_irqc =
      (
         ({CONFIG_DW{msr_irqc_imr_sel}} & msr_irqc_imr) |
         ({CONFIG_DW{msr_irqc_irr_sel}} & msr_irqc_irr)
      );
   assign msr_tsc_tsr_sel = s1i_bank_off[0];
   assign msr_tsc_tcr_sel = s1i_bank_off[1];
   assign dout_tsc =
      (
         ({CONFIG_DW{msr_tsc_tsr_sel}} & msr_tsc_tsr) |
         ({CONFIG_DW{msr_tsc_tcr_sel}} & msr_tsc_tcr)
      );
   ysyx_20210479_pmux #(.SELW(4), .DW(CONFIG_DW)) pmux_dout_sr (.sel(s1i_bank_off[4-1:0]), .din(msr_sr), .dout(dout_sr));
   assign s1i_bank_ps = (s1i_bank_addr == 0);
   assign s1i_bank_imm = (s1i_bank_addr == 1);
   assign s1i_bank_dmm = (s1i_bank_addr == 2);
   assign s1i_bank_ic = (s1i_bank_addr == 3);
   assign s1i_bank_dc = (s1i_bank_addr == 4);
   assign s1i_bank_dbg = (s1i_bank_addr == 5);
   assign s1i_bank_irqc = (s1i_bank_addr == 6);
   assign s1i_bank_tsc = (s1i_bank_addr == 7);
   assign s1i_bank_sr = (s1i_bank_addr == 8);
   assign epu_dout =
      (
         ({CONFIG_DW{s1i_bank_ps}} & dout_ps) |
         ({CONFIG_DW{s1i_bank_imm}} & dout_imm) |
         ({CONFIG_DW{s1i_bank_dmm}} & dout_dmm) |
         ({CONFIG_DW{s1i_bank_ic}} & dout_ic) |
         ({CONFIG_DW{s1i_bank_dc}} & dout_dc) |
         ({CONFIG_DW{s1i_bank_irqc}} & dout_irqc) |
         ({CONFIG_DW{s1i_bank_tsc}} & dout_tsc) |
         ({CONFIG_DW{s1i_bank_sr}} & dout_sr)
      );
   assign epu_dout_valid = (ex_valid & ~flush_s1 & ex_epu_opc_bus[1]);
   assign s1i_ERET = (ex_valid & ~flush_s1 & ex_epu_opc_bus[3]);
   assign s1i_ESYSCALL = (ex_valid & ~flush_s1 & ex_epu_opc_bus[2]);
   assign s1i_EINSN = (ex_valid & ~flush_s1 & ex_epu_opc_bus[(8-1)]);
   assign s1i_EIPF = (ex_valid & ~flush_s1 & ex_epu_opc_bus[5]);
   assign s1i_EITM = (ex_valid & ~flush_s1 & ex_epu_opc_bus[4]);
   assign s1i_EIRQ = (ex_valid & ~flush_s1 & ex_epu_opc_bus[6]);
   assign s1i_E_FLUSH_TLB = (ex_valid & ~flush_s1 & (s1i_wmsr_psr_we |
                              s1i_msr_imm_tlbl_we |
                              s1i_msr_imm_tlbh_we |
                              s1i_msr_dmm_tlbl_we |
                              s1i_msr_dmm_tlbh_we));
   assign s1i_wmsr_psr_we      = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_ps & s1i_bank_off[0];
   assign s1i_wmsr_epc_we      = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_ps & s1i_bank_off[3];
   assign s1i_wmsr_epsr_we     = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_ps & s1i_bank_off[2];
   assign s1i_wmsr_elsa_we     = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_ps & s1i_bank_off[4];
   assign s1i_msr_imm_tlbl_we  = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_imm & msr_imm_tlbl_sel;
   assign s1i_msr_imm_tlbh_we  = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_imm & msr_imm_tlbh_sel;
   assign s1i_msr_dmm_tlbl_we  = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_dmm & msr_dmm_tlbl_sel;
   assign s1i_msr_dmm_tlbh_we  = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_dmm & msr_dmm_tlbh_sel;
   assign s1i_msr_ic_inv_we    = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_ic & msr_ic_inv_sel;
   assign s1i_msr_dc_inv_we    = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_dc & msr_dc_inv_sel;
   assign s1i_msr_dc_fls_we    = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_dc & msr_dc_fls_sel;
   assign s1i_msr_irqc_imr_we  = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_irqc & msr_irqc_imr_sel;
   assign s1i_msr_tsc_tsr_we   = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_tsc & msr_tsc_tsr_sel;
   assign s1i_msr_tsc_tcr_we   = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_tsc & msr_tsc_tcr_sel;
   assign s1i_msr_sr_we        = ex_valid & ~flush_s1 & ex_epu_opc_bus[0] & s1i_bank_sr;
   assign s1i_wmsr_we = {s1i_wmsr_psr_we,
                        s1i_wmsr_epc_we,
                        s1i_wmsr_epsr_we,
                        s1i_wmsr_elsa_we,
                        s1i_msr_imm_tlbl_we,
                        s1i_msr_imm_tlbh_we,
                        s1i_msr_dmm_tlbl_we,
                        s1i_msr_dmm_tlbh_we,
                        s1i_msr_irqc_imr_we,
                        s1i_msr_tsc_tsr_we,
                        s1i_msr_tsc_tcr_we,
                        s1i_msr_sr_we,
                        s1i_bank_off};
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_ERET (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_ERET), .Q(s1o_commit_ERET) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_ESYSCALL (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_ESYSCALL), .Q(s1o_commit_ESYSCALL) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_EINSN (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_EINSN), .Q(s1o_commit_EINSN) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_EIPF (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_EIPF), .Q(s1o_commit_EIPF) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_EITM (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_EITM), .Q(s1o_commit_EITM) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_EIRQ (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_EIRQ), .Q(s1o_commit_EIRQ) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_commit_E_FLUSH_TLB (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_E_FLUSH_TLB), .Q(s1o_commit_E_FLUSH_TLB) );
   ysyx_20210479_mDFF_lr # (.DW(NCPU_WMSR_WE_W)) ff_s1o_commit_wmsr_we (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_wmsr_we), .Q(s1o_commit_wmsr_we) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW)) ff_s1o_commit_wmsr_dat (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_msr_wdat), .Q(s1o_commit_wmsr_dat) );
   ysyx_20210479_mDFF_l # (.DW((CONFIG_AW-2 ))) ff_s1o_commit_epc (.CLK(clk), .LOAD(p_ce_s1), .D(ex_pc), .Q(s1o_commit_epc) );
   ysyx_20210479_mDFF_l # (.DW((CONFIG_AW-2 ))) ff_s1o_commit_nepc (.CLK(clk), .LOAD(p_ce_s1), .D(ex_npc), .Q(s1o_commit_nepc) );
   assign {
      s1o_commit_wmsr_psr_we,
      s1o_commit_wmsr_epc_we,
      s1o_commit_wmsr_epsr_we,
      s1o_commit_wmsr_elsa_we,
      s1o_commit_msr_imm_tlbl_we,
      s1o_commit_msr_imm_tlbh_we,
      s1o_commit_msr_dmm_tlbl_we,
      s1o_commit_msr_dmm_tlbh_we,
      s1o_commit_msr_irqc_imr_we,
      s1o_commit_msr_tsc_tsr_we,
      s1o_commit_msr_tsc_tcr_we,
      s1o_commit_msr_sr_we,
      s1o_commit_bank_off} = ({NCPU_WMSR_WE_W{p_ce_s2}} & s1o_commit_wmsr_we);
   assign {s1o_wmsr_psr_dce,s1o_wmsr_psr_ice,s1o_wmsr_psr_dmme,s1o_wmsr_psr_imme,s1o_wmsr_psr_ire,s1o_wmsr_psr_rm} = s1o_commit_wmsr_dat[9:4];
   assign msr_psr_save = (p_ce_s2 & (s1o_commit_ESYSCALL |
                                    s1o_commit_EITM |
                                    s1o_commit_EIPF |
                                    s1o_commit_EINSN |
                                    s2i_EDTM |
                                    s2i_EDPF |
                                    s2i_EALIGN |
                                    s1o_commit_EIRQ));
   assign msr_psr_restore = (p_ce_s2 & s1o_commit_ERET);
   assign msr_psr_rm_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_rm_nxt = s1o_wmsr_psr_rm;
   assign msr_psr_imme_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_imme_nxt = s1o_wmsr_psr_imme;
   assign msr_psr_dmme_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_dmme_nxt = s1o_wmsr_psr_dmme;
   assign msr_psr_ire_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_ire_nxt = s1o_wmsr_psr_ire;
   assign msr_psr_ice_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_ice_nxt = s1o_wmsr_psr_ice;
   assign msr_psr_dce_we = s1o_commit_wmsr_psr_we;
   assign msr_psr_dce_nxt = s1o_wmsr_psr_dce;
   assign msr_epsr_we = s1o_commit_wmsr_epsr_we;
   assign msr_epsr_nxt = s1o_commit_wmsr_dat[10-1:0];
   assign msr_epc_nxt = (s1o_commit_wmsr_epc_we)
                           ? s1o_commit_wmsr_dat
                           : (s1o_commit_ESYSCALL)
                              ? {s1o_commit_nepc,2'b0}
                              : {s1o_commit_epc,2'b0};
   assign msr_epc_we = (msr_psr_save | s1o_commit_wmsr_epc_we);
   assign s1o_set_elsa_as_pc = (s1o_commit_EITM | s1o_commit_EIPF | s1o_commit_EINSN);
   assign s1o_set_elsa = (s1o_set_elsa_as_pc | s2i_EDTM | s2i_EDPF | s2i_EALIGN);
   assign s1o_lsa_nxt = s1o_set_elsa_as_pc ? {s1o_commit_epc,2'b0} : s2i_vaddr;
   assign msr_elsa_nxt = s1o_set_elsa ? s1o_lsa_nxt : s1o_commit_wmsr_dat;
   assign msr_elsa_we = s1o_set_elsa | s1o_commit_wmsr_elsa_we;
   assign msr_imm_tlbl_idx = s1o_commit_bank_off[CONFIG_ITLB_P_SETS-1:0];
   assign msr_imm_tlbl_nxt = s1o_commit_wmsr_dat;
   assign msr_imm_tlbl_we = s1o_commit_msr_imm_tlbl_we;
   assign msr_imm_tlbh_idx = s1o_commit_bank_off[CONFIG_ITLB_P_SETS-1:0];
   assign msr_imm_tlbh_nxt = s1o_commit_wmsr_dat;
   assign msr_imm_tlbh_we = s1o_commit_msr_imm_tlbh_we;
   assign msr_dmm_tlbl_idx = s1o_commit_bank_off[CONFIG_DTLB_P_SETS-1:0];
   assign msr_dmm_tlbl_nxt = s1o_commit_wmsr_dat;
   assign msr_dmm_tlbl_we = s1o_commit_msr_dmm_tlbl_we;
   assign msr_dmm_tlbh_idx = s1o_commit_bank_off[CONFIG_DTLB_P_SETS-1:0];
   assign msr_dmm_tlbh_nxt = s1o_commit_wmsr_dat;
   assign msr_dmm_tlbh_we = s1o_commit_msr_dmm_tlbh_we;
   assign msr_icinv_we = (s1i_msr_ic_inv_we & p_ce_s1_no_icinv_stall);
   assign msr_icinv_nxt = s1i_msr_wdat;
   assign msr_dcinv_we = s1i_msr_dc_inv_we;
   assign msr_dcinv_nxt = s1i_msr_wdat;
   assign msr_dcfls_we = s1i_msr_dc_fls_we;
   assign msr_dcfls_nxt = s1i_msr_wdat;
   assign msr_irqc_imr_we = s1o_commit_msr_irqc_imr_we;
   assign msr_irqc_imr_nxt = s1o_commit_wmsr_dat;
   assign msr_tsc_tsr_we = s1o_commit_msr_tsc_tsr_we;
   assign msr_tsc_tsr_nxt = s1o_commit_wmsr_dat;
   assign msr_tsc_tcr_we = s1o_commit_msr_tsc_tcr_we;
   assign msr_tsc_tcr_nxt = s1o_commit_wmsr_dat;
   assign msr_sr_we = (s1o_commit_bank_off[4-1:0] & {4{s1o_commit_msr_sr_we}});
   assign msr_sr_nxt = s1o_commit_wmsr_dat;
   assign exc_flush_tgt = ({(CONFIG_AW-2 ){s2i_EDTM}} & CONFIG_EDTM_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s2i_EDPF}} & CONFIG_EDPF_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s2i_EALIGN}} & CONFIG_EALIGN_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_E_FLUSH_TLB}} & s1o_commit_nepc) |
                           ({(CONFIG_AW-2 ){s1o_commit_ESYSCALL}} & CONFIG_ESYSCALL_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_ERET}} & msr_epc[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_EITM}} & CONFIG_EITM_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_EIPF}} & CONFIG_EIPF_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_EIRQ}} & CONFIG_EIRQ_VECTOR[2  +: (CONFIG_AW-2 )]) |
                           ({(CONFIG_AW-2 ){s1o_commit_EINSN}} & CONFIG_EINSN_VECTOR[2  +: (CONFIG_AW-2 )]);
   assign exc_flush = p_ce_s2 & (s2i_EDTM |
                        s2i_EDPF |
                        s2i_EALIGN |
                        s1o_commit_E_FLUSH_TLB |
                        s1o_commit_ESYSCALL |
                        s1o_commit_ERET |
                        s1o_commit_EITM |
                        s1o_commit_EIPF |
                        s1o_commit_EIRQ |
                        s1o_commit_EINSN);
   ysyx_20210479_ex_epu_irqc
      #(
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_NUM_IRQ                 (CONFIG_NUM_IRQ))
   U_IRQC
      (
       .irq_async                       (irq_async),
       .msr_irqc_imr                    (msr_irqc_imr[CONFIG_DW-1:0]),
       .msr_irqc_irr                    (msr_irqc_irr[CONFIG_DW-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .irqs                            (irqs[CONFIG_NUM_IRQ-1:0]),
       .msr_psr_ire                     (msr_psr_ire),
       .msr_irqc_imr_nxt                (msr_irqc_imr_nxt[CONFIG_DW-1:0]),
       .msr_irqc_imr_we                 (msr_irqc_imr_we));
   ysyx_20210479_ex_epu_tsc
      #(
        .CONFIG_DW                      (CONFIG_DW))
   U_TSC
      (
       .tsc_irq                         (tsc_irq),
       .msr_tsc_tsr                     (msr_tsc_tsr[CONFIG_DW-1:0]),
       .msr_tsc_tcr                     (msr_tsc_tcr[CONFIG_DW-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .msr_tsc_tsr_nxt                 (msr_tsc_tsr_nxt[CONFIG_DW-1:0]),
       .msr_tsc_tsr_we                  (msr_tsc_tsr_we),
       .msr_tsc_tcr_nxt                 (msr_tsc_tcr_nxt[CONFIG_DW-1:0]),
       .msr_tsc_tcr_we                  (msr_tsc_tcr_we));
endmodule
module ysyx_20210479_ex_epu_irqc
#(
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_NUM_IRQ = 0
)
(
   input                               clk,
   input                               rst,
   input [CONFIG_NUM_IRQ-1:0]          irqs,
   output                              irq_async,
   input                               msr_psr_ire,
   output [CONFIG_DW-1:0]              msr_irqc_imr,
   input [CONFIG_DW-1:0]               msr_irqc_imr_nxt,
   input                               msr_irqc_imr_we,
   output [CONFIG_DW-1:0]              msr_irqc_irr
);
   wire [CONFIG_DW-1:0]                imr_ff;
   wire [CONFIG_NUM_IRQ-1:0]           msr_irqc_irr_0;
   wire [CONFIG_NUM_IRQ-1:0]           irq_masked;
   ysyx_20210479_mDFF_r #(CONFIG_NUM_IRQ) dff_msr_irqc_irr_0 (.CLK(clk), .RST(rst), .D(irqs), .Q(msr_irqc_irr_0) );
   ysyx_20210479_mDFF_r #(CONFIG_NUM_IRQ) dff_msr_irqc_irr (.CLK(clk), .RST(rst), .D(msr_irqc_irr_0), .Q(msr_irqc_irr) );
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_DW), .RST_VECTOR({CONFIG_DW{1'b1}})) ff_imr_ (.CLK(clk), .RST(rst), .LOAD(msr_irqc_imr_we), .D(msr_irqc_imr_nxt), .Q(imr_ff) );
   assign msr_irqc_imr = (msr_irqc_imr_we) ? msr_irqc_imr_nxt : imr_ff;
   assign irq_masked = (msr_irqc_irr & ~msr_irqc_imr);
   assign irq_async = (|irq_masked & msr_psr_ire);
endmodule
module ysyx_20210479_ex_epu_tsc
#(
   parameter                           CONFIG_DW = 0
)
(
   input                               clk,
   input                               rst,
   output                              tsc_irq,
   output [CONFIG_DW-1:0]              msr_tsc_tsr,
   input [CONFIG_DW-1:0]               msr_tsc_tsr_nxt,
   input                               msr_tsc_tsr_we,
   output [CONFIG_DW-1:0]              msr_tsc_tcr,
   input [CONFIG_DW-1:0]               msr_tsc_tcr_nxt,
   input                               msr_tsc_tcr_we
);
   wire [CONFIG_DW-1:0]                tcr_ff;
   wire [CONFIG_DW-1:0]                msr_tsc_tcr_ff;
   wire [28-1:0]         tcr_cnt;
   wire                                tcr_en;
   wire                                tcr_i;
   wire                                tcr_p;
   wire                                count;
   wire                                count_clk;
   wire [CONFIG_DW-1:0]                tsr_nxt;
   wire                                irq_set;
   wire                                irq_clr;
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_DW)) ff_tcr (.CLK(clk), .RST(rst), .LOAD(msr_tsc_tcr_we), .D(msr_tsc_tcr_nxt), .Q(tcr_ff) );
   assign msr_tsc_tcr_ff[28-1:0] = tcr_ff[28-1:0];
   assign msr_tsc_tcr_ff[28] = tcr_ff[28];
   assign msr_tsc_tcr_ff[29] = tcr_ff[29];
   assign msr_tsc_tcr_ff[30] = tsc_irq;
   assign msr_tsc_tcr_ff[31] = tcr_ff[31];
   assign msr_tsc_tcr = msr_tsc_tcr_we ? msr_tsc_tcr_nxt : msr_tsc_tcr_ff;
   assign tcr_cnt = msr_tsc_tcr[28-1:0];
   assign tcr_en = msr_tsc_tcr[28];
   assign tcr_i = msr_tsc_tcr[29];
   assign tcr_p = msr_tsc_tcr[30];
   assign count = tcr_en;
   assign count_clk = clk;
   assign tsr_nxt = msr_tsc_tsr_we ? msr_tsc_tsr_nxt : msr_tsc_tsr+1'b1;
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_DW)) ff_msr_tsc_tsr (.CLK(count_clk), .RST(rst), .LOAD(msr_tsc_tsr_we|count), .D(tsr_nxt), .Q(msr_tsc_tsr) );
   assign irq_set = (msr_tsc_tsr[28-1:0]==tcr_cnt) & tcr_i;
   assign irq_clr = msr_tsc_tcr_we & ~tcr_p;
   ysyx_20210479_mDFF_lr #(1) ff_tsc_irq (.CLK(clk), .RST(rst), .LOAD(irq_set|irq_clr), .D(irq_set & ~irq_clr), .Q(tsc_irq) );
endmodule
module ysyx_20210479_ex_lsu
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_DW = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_DMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_DTLB_P_SETS = 0,
   parameter                           CONFIG_DC_P_LINE = 0,
   parameter                           CONFIG_DC_P_SETS = 0,
   parameter                           CONFIG_DC_P_WAYS = 0,
   parameter                           AXI_P_DW_BYTES    = 0,
   parameter                           AXI_ADDR_WIDTH    = 0,
   parameter                           AXI_ID_WIDTH      = 0,
   parameter                           AXI_USER_WIDTH    = 0
)
(
   input                               clk,
   input                               rst,
   input                               p_ce_s1,
   input                               flush_s1,
   output                              lsu_stall_req,
   input                               ex_valid,
   input [7-1:0]          ex_lsu_opc_bus,
   output                              agu_en,
   input [CONFIG_DW-1:0]               add_sum,
   input [CONFIG_DW-1:0]               ex_operand2,
   input                               dbus_ARREADY,
   output                              dbus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_ARADDR,
   output [2:0]                        dbus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_ARID,
   output [AXI_USER_WIDTH-1:0]         dbus_ARUSER,
   output [7:0]                        dbus_ARLEN,
   output [2:0]                        dbus_ARSIZE,
   output [1:0]                        dbus_ARBURST,
   output                              dbus_ARLOCK,
   output [3:0]                        dbus_ARCACHE,
   output [3:0]                        dbus_ARQOS,
   output [3:0]                        dbus_ARREGION,
   output                              dbus_RREADY,
   input                               dbus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_RDATA,
   input  [1:0]                        dbus_RRESP,
   input                               dbus_RLAST,
   input  [AXI_ID_WIDTH-1:0]           dbus_RID,
   input  [AXI_USER_WIDTH-1:0]         dbus_RUSER,
   input                               dbus_AWREADY,
   output                              dbus_AWVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_AWADDR,
   output [2:0]                        dbus_AWPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_AWID,
   output [AXI_USER_WIDTH-1:0]         dbus_AWUSER,
   output [7:0]                        dbus_AWLEN,
   output [2:0]                        dbus_AWSIZE,
   output [1:0]                        dbus_AWBURST,
   output                              dbus_AWLOCK,
   output [3:0]                        dbus_AWCACHE,
   output [3:0]                        dbus_AWQOS,
   output [3:0]                        dbus_AWREGION,
   input                               dbus_WREADY,
   output                              dbus_WVALID,
   output [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_WDATA,
   output [(1<<AXI_P_DW_BYTES)-1:0]    dbus_WSTRB,
   output                              dbus_WLAST,
   output [AXI_USER_WIDTH-1:0]         dbus_WUSER,
   output                              dbus_BREADY,
   input                               dbus_BVALID,
   input [1:0]                         dbus_BRESP,
   input [AXI_ID_WIDTH-1:0]            dbus_BID,
   input [AXI_USER_WIDTH-1:0]          dbus_BUSER,
   output                              lsu_EDTM,
   output                              lsu_EDPF,
   output                              lsu_EALIGN,
   output [CONFIG_AW-1:0]              lsu_vaddr,
   output [CONFIG_DW-1:0]              lsu_dout,
   input                               msr_psr_dmme,
   input                               msr_psr_rm,
   input                               msr_psr_dce,
   output [CONFIG_DW-1:0]              msr_dmmid,
   input [CONFIG_DTLB_P_SETS-1:0]      msr_dmm_tlbl_idx,
   input [CONFIG_DW-1:0]               msr_dmm_tlbl_nxt,
   input                               msr_dmm_tlbl_we,
   input [CONFIG_DTLB_P_SETS-1:0]      msr_dmm_tlbh_idx,
   input [CONFIG_DW-1:0]               msr_dmm_tlbh_nxt,
   input                               msr_dmm_tlbh_we,
   output [CONFIG_DW-1:0]              msr_dcid,
   input [CONFIG_DW-1:0]               msr_dcinv_nxt,
   input                               msr_dcinv_we,
   input [CONFIG_DW-1:0]               msr_dcfls_nxt,
   input                               msr_dcfls_we
);
   localparam CONFIG_P_DW_BYTES        = (CONFIG_P_DW-3);
   wire                 dc_stall_req;           
   wire                                s1i_valid;
   wire                                s1i_load;
   wire                                s1i_store;
   wire                                s1i_sign_ext;
   wire                                s1i_barr;
   wire                                s1i_dcop;
   wire                                s1i_dc_req;
   wire                                s1i_tlb_req;
   wire [CONFIG_AW-1:0]                s1i_dc_vaddr;
   wire [CONFIG_P_PAGE_SIZE-1:0]       s1i_dc_vpo;
   wire [CONFIG_DW/8-1:0]              s1i_dc_wmsk;
   wire [CONFIG_DW-1:0]                s1i_dc_wdat;
   wire                                s1i_misalign;
   wire [CONFIG_DW-1:0]                s1i_din_8b;
   wire [CONFIG_DW-1:0]                s1i_din_16b;
   wire [3:0]                          s1i_we_msk_8b;
   wire [3:0]                          s1i_we_msk_16b;
   wire [2:0]                          s1i_size;
   wire                                s1o_valid;
   wire [2:0]                          s1o_size;
   wire                                s1o_sign_ext;
   wire                                s2i_tlb_uncached;
   wire                                s2i_tlb_exc;
   wire                                s2i_kill_req;
   wire                                s2i_uncached;
   wire [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] s2i_tlb_ppn;
   wire [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] s2i_dc_ppn;
   wire                                s1o_EDTM;
   wire                                s1o_EDPF;
   wire                                s1o_EALIGN;
   wire [CONFIG_AW-1:0]                s1o_vaddr;
   wire                                s1o_dcop;
   wire                                s1o_msr_psr_dce;
   wire [CONFIG_DW-1:0]                s2o_dout_32b;
   wire [7:0]                          s2o_dout_8b;
   wire [15:0]                         s2o_dout_16b;
   wire [CONFIG_AW-1:0]                s2o_vaddr;
   wire [2:0]                          s2o_size;
   wire                                s2o_sign_ext;
   assign s1i_valid = ex_valid & ~flush_s1 & (s1i_load|s1i_store|s1i_dcop);
   assign s1i_load = ex_lsu_opc_bus[0];
   assign s1i_store = ex_lsu_opc_bus[1];
   assign s1i_sign_ext = ex_lsu_opc_bus[3];
   assign s1i_barr = ex_lsu_opc_bus[2];
   assign s1i_size = ex_lsu_opc_bus[6:4];
   assign s1i_dcop = (msr_dcinv_we | msr_dcfls_we);
   assign agu_en = (s1i_load|s1i_store);
   assign s1i_dc_vaddr = (msr_dcinv_we)
                           ? msr_dcinv_nxt
                           : (msr_dcfls_we)
                              ? msr_dcfls_nxt
                              : add_sum;
   assign s1i_misalign = (s1i_size==3'd3 & |s1i_dc_vaddr[1:0]) |
                           (s1i_size==3'd2 & s1i_dc_vaddr[0]);
   assign s1i_din_8b = {ex_operand2[7:0], ex_operand2[7:0], ex_operand2[7:0], ex_operand2[7:0]};
   assign s1i_din_16b = {ex_operand2[15:0], ex_operand2[15:0]};
   assign s1i_dc_wdat = ({CONFIG_DW{s1i_size==3'd3}} & ex_operand2) |
                        ({CONFIG_DW{s1i_size==3'd2}} & s1i_din_16b) |
                        ({CONFIG_DW{s1i_size==3'd1}} & s1i_din_8b);
   assign s1i_we_msk_8b = (s1i_dc_vaddr[1:0]==2'b00 ? 4'b0001 :
                           s1i_dc_vaddr[1:0]==2'b01 ? 4'b0010 :
                           s1i_dc_vaddr[1:0]==2'b10 ? 4'b0100 :
                           s1i_dc_vaddr[1:0]==2'b11 ? 4'b1000 : 4'b0000);
   assign s1i_we_msk_16b = s1i_dc_vaddr[1] ? 4'b1100 : 4'b0011;
   assign s1i_dc_wmsk = {CONFIG_DW/8{s1i_store}} & (
                        ({CONFIG_DW/8{s1i_size==3'd3}} & 4'b1111) |
                        ({CONFIG_DW/8{s1i_size==3'd2}} & s1i_we_msk_16b) |
                        ({CONFIG_DW/8{s1i_size==3'd1}} & s1i_we_msk_8b) );
   assign s1i_dc_vpo = s1i_dc_vaddr[CONFIG_P_PAGE_SIZE-1:0];
   assign s1i_dc_req = (p_ce_s1 & s1i_valid);
   assign s1i_tlb_req = (s1i_dc_req & ~s1i_dcop);
   ysyx_20210479_dmmu
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_DMMU_ENABLE_UNCACHED_SEG(CONFIG_DMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_DTLB_P_SETS             (CONFIG_DTLB_P_SETS))
   U_D_MMU
      (
         .clk                          (clk),
         .rst                          (rst),
         .re                           (s1i_tlb_req),
         .vpn                          (s1i_dc_vaddr[CONFIG_AW-1:CONFIG_P_PAGE_SIZE]),
         .we                           (s1i_store),
         .ppn                          (s2i_tlb_ppn),
         .EDTM                         (s1o_EDTM),
         .EDPF                         (s1o_EDPF),
         .uncached                     (s2i_tlb_uncached),
         .msr_psr_dmme                 (msr_psr_dmme),
         .msr_psr_rm                   (msr_psr_rm),
         .msr_dmmid                    (msr_dmmid),
         .msr_dmm_tlbl_idx             (msr_dmm_tlbl_idx),
         .msr_dmm_tlbl_nxt             (msr_dmm_tlbl_nxt),
         .msr_dmm_tlbl_we              (msr_dmm_tlbl_we),
         .msr_dmm_tlbh_idx             (msr_dmm_tlbh_idx),
         .msr_dmm_tlbh_nxt             (msr_dmm_tlbh_nxt),
         .msr_dmm_tlbh_we              (msr_dmm_tlbh_we)
      );
   assign s2i_tlb_exc = (s1o_EDTM | s1o_EDPF | s1o_EALIGN);
   assign s2i_kill_req = (s2i_tlb_exc);
   assign s2i_uncached = (s2i_tlb_uncached | ~s1o_msr_psr_dce);
   assign s2i_dc_ppn = (s1o_dcop)
                        ? s1o_vaddr[CONFIG_AW-1:CONFIG_P_PAGE_SIZE]
                        : s2i_tlb_ppn;
   ysyx_20210479_dcache
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_DW                    (CONFIG_P_DW),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_DC_P_LINE               (CONFIG_DC_P_LINE),
        .CONFIG_DC_P_SETS               (CONFIG_DC_P_SETS),
        .CONFIG_DC_P_WAYS               (CONFIG_DC_P_WAYS),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_D_CACHE
      (
       .stall_req                       (dc_stall_req),          
       .dout                            (s2o_dout_32b),          
       .dbus_ARVALID                    (dbus_ARVALID),
       .dbus_ARADDR                     (dbus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_ARPROT                     (dbus_ARPROT[2:0]),
       .dbus_ARID                       (dbus_ARID[AXI_ID_WIDTH-1:0]),
       .dbus_ARUSER                     (dbus_ARUSER[AXI_USER_WIDTH-1:0]),
       .dbus_ARLEN                      (dbus_ARLEN[7:0]),
       .dbus_ARSIZE                     (dbus_ARSIZE[2:0]),
       .dbus_ARBURST                    (dbus_ARBURST[1:0]),
       .dbus_ARLOCK                     (dbus_ARLOCK),
       .dbus_ARCACHE                    (dbus_ARCACHE[3:0]),
       .dbus_ARQOS                      (dbus_ARQOS[3:0]),
       .dbus_ARREGION                   (dbus_ARREGION[3:0]),
       .dbus_RREADY                     (dbus_RREADY),
       .dbus_AWVALID                    (dbus_AWVALID),
       .dbus_AWADDR                     (dbus_AWADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_AWPROT                     (dbus_AWPROT[2:0]),
       .dbus_AWID                       (dbus_AWID[AXI_ID_WIDTH-1:0]),
       .dbus_AWUSER                     (dbus_AWUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWLEN                      (dbus_AWLEN[7:0]),
       .dbus_AWSIZE                     (dbus_AWSIZE[2:0]),
       .dbus_AWBURST                    (dbus_AWBURST[1:0]),
       .dbus_AWLOCK                     (dbus_AWLOCK),
       .dbus_AWCACHE                    (dbus_AWCACHE[3:0]),
       .dbus_AWQOS                      (dbus_AWQOS[3:0]),
       .dbus_AWREGION                   (dbus_AWREGION[3:0]),
       .dbus_WVALID                     (dbus_WVALID),
       .dbus_WDATA                      (dbus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_WSTRB                      (dbus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]),
       .dbus_WLAST                      (dbus_WLAST),
       .dbus_WUSER                      (dbus_WUSER[AXI_USER_WIDTH-1:0]),
       .dbus_BREADY                     (dbus_BREADY),
       .msr_dcid                        (msr_dcid[CONFIG_DW-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .req                             (s1i_dc_req),            
       .size                            (s1i_size),              
       .wmsk                            (s1i_dc_wmsk),           
       .wdat                            (s1i_dc_wdat),           
       .vpo                             (s1i_dc_vpo),            
       .ppn_s2                          (s2i_dc_ppn),            
       .kill_req_s2                     (s2i_kill_req),          
       .uncached_s2                     (s2i_uncached),          
       .inv                             (msr_dcinv_we),          
       .fls                             (msr_dcfls_we),          
       .dbus_ARREADY                    (dbus_ARREADY),
       .dbus_RVALID                     (dbus_RVALID),
       .dbus_RDATA                      (dbus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_RLAST                      (dbus_RLAST),
       .dbus_AWREADY                    (dbus_AWREADY),
       .dbus_WREADY                     (dbus_WREADY),
       .dbus_BVALID                     (dbus_BVALID),
       .dbus_RRESP                      (dbus_RRESP[1:0]),
       .dbus_RID                        (dbus_RID[AXI_ID_WIDTH-1:0]),
       .dbus_RUSER                      (dbus_RUSER[AXI_USER_WIDTH-1:0]),
       .dbus_BRESP                      (dbus_BRESP[1:0]),
       .dbus_BID                        (dbus_BID[AXI_ID_WIDTH-1:0]),
       .dbus_BUSER                      (dbus_BUSER[AXI_USER_WIDTH-1:0]));
   ysyx_20210479_mDFF_l #(.DW(3)) ff_s1o_size (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_size), .Q(s1o_size) );
   ysyx_20210479_mDFF_l #(.DW(CONFIG_AW)) ff_s1o_vaddr (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_dc_vaddr), .Q(s1o_vaddr) );
   ysyx_20210479_mDFF_l #(.DW(1)) ff_s1o_sign_ext (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_sign_ext), .Q(s1o_sign_ext) );
   ysyx_20210479_mDFF_l #(.DW(1)) ff_s1o_dcop (.CLK(clk), .LOAD(p_ce_s1), .D(s1i_dcop), .Q(s1o_dcop) );
   ysyx_20210479_mDFF_l #(.DW(CONFIG_AW)) ff_s2o_vaddr (.CLK(clk), .LOAD(p_ce_s1), .D(s1o_vaddr), .Q(s2o_vaddr) );
   ysyx_20210479_mDFF_l #(.DW(3)) ff_s2o_size (.CLK(clk), .LOAD(p_ce_s1), .D(s1o_size), .Q(s2o_size) );
   ysyx_20210479_mDFF_l #(.DW(1)) ff_s2o_sign_ext (.CLK(clk), .LOAD(p_ce_s1), .D(s1o_sign_ext), .Q(s2o_sign_ext) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_s1o_valid (.CLK(clk), .RST(rst), .LOAD(p_ce_s1|flush_s1), .D(s1i_valid), .Q(s1o_valid) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_s1o_misalign (.CLK(clk), .RST(rst), .LOAD(p_ce_s1), .D(s1i_misalign), .Q(s1o_EALIGN) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_s1o_msr_psr_dce (.CLK(clk), .RST(rst), .LOAD(p_ce_s1), .D(msr_psr_dce), .Q(s1o_msr_psr_dce) );
   assign lsu_stall_req = (dc_stall_req);
   assign s2o_dout_8b = ({8{s2o_vaddr[1:0]==2'b00}} & s2o_dout_32b[7:0]) |
                          ({8{s2o_vaddr[1:0]==2'b01}} & s2o_dout_32b[15:8]) |
                          ({8{s2o_vaddr[1:0]==2'b10}} & s2o_dout_32b[23:16]) |
                          ({8{s2o_vaddr[1:0]==2'b11}} & s2o_dout_32b[31:24]);
   assign s2o_dout_16b = s2o_vaddr[1] ? s2o_dout_32b[31:16] : s2o_dout_32b[15:0];
   assign lsu_dout =
      ({CONFIG_DW{s2o_size==3'd3}} & s2o_dout_32b) |
      ({CONFIG_DW{s2o_size==3'd2}} & {{16{s2o_sign_ext & s2o_dout_16b[15]}}, s2o_dout_16b[15:0]}) |
      ({CONFIG_DW{s2o_size==3'd1}} & {{24{s2o_sign_ext & s2o_dout_8b[7]}}, s2o_dout_8b[7:0]});
   assign lsu_EDTM = (s1o_valid & s1o_EDTM);
   assign lsu_EDPF = (s1o_valid & s1o_EDPF);
   assign lsu_EALIGN = (s1o_valid & s1o_EALIGN);
   assign lsu_vaddr = s1o_vaddr;
endmodule
module ysyx_20210479_ex_psr
#(
   parameter                           CONFIG_DW = 0,
   parameter [7:0]                     CPUID_VER = 1,
   parameter [9:0]                     CPUID_REV = 0,
   parameter [0:0]                     CPUID_FIMM = 1,
   parameter [0:0]                     CPUID_FDMM = 1,
   parameter [0:0]                     CPUID_FICA = 0,
   parameter [0:0]                     CPUID_FDCA = 0,
   parameter [0:0]                     CPUID_FDBG = 0,
   parameter [0:0]                     CPUID_FFPU = 0,
   parameter [0:0]                     CPUID_FIRQC = 1,
   parameter [0:0]                     CPUID_FTSC = 1
)
(
   input                               clk,
   input                               rst,
   input                               msr_psr_save,
   input                               msr_psr_restore,
   output [10-1:0]           msr_psr,
   input                               msr_psr_rm_nxt,
   output                              msr_psr_rm,
   input                               msr_psr_rm_we,
   input                               msr_psr_ire_nxt,
   output                              msr_psr_ire,
   input                               msr_psr_ire_we,
   input                               msr_psr_imme_nxt,
   output                              msr_psr_imme,
   input                               msr_psr_imme_we,
   input                               msr_psr_dmme_nxt,
   output                              msr_psr_dmme,
   input                               msr_psr_dmme_we,
   input                               msr_psr_ice_nxt,
   output                              msr_psr_ice,
   input                               msr_psr_ice_we,
   input                               msr_psr_dce_nxt,
   output                              msr_psr_dce,
   input                               msr_psr_dce_we,
   output [CONFIG_DW-1:0]              msr_cpuid,
   input [10-1:0]            msr_epsr_nxt,
   output [10-1:0]           msr_epsr,
   input                               msr_epsr_we,
   input [CONFIG_DW-1:0]               msr_epc_nxt,
   output [CONFIG_DW-1:0]              msr_epc,
   input                               msr_epc_we,
   input [CONFIG_DW-1:0]               msr_elsa_nxt,
   output [CONFIG_DW-1:0]              msr_elsa,
   input                               msr_elsa_we,
   output [CONFIG_DW-1:0]              msr_coreid,
   output [CONFIG_DW*4-1:0] msr_sr,
   input [CONFIG_DW-1:0]               msr_sr_nxt,
   input [4-1:0]            msr_sr_we
);
   wire                                msr_psr_rm_ff;
   wire                                msr_psr_ire_ff;
   wire                                msr_psr_imme_ff;
   wire                                msr_psr_dmme_ff;
   wire                                msr_psr_rm_nold;
   wire                                msr_psr_ire_nold;
   wire                                msr_psr_imme_nold;
   wire                                msr_psr_dmme_nold;
   wire                                msr_psr_ice_ff;
   wire                                msr_psr_dce_ff;
   wire [10-1:0]             msr_psr_nold;
   wire [10-1:0]             msr_epsr_ff;
   wire [CONFIG_DW-1:0]                msr_epc_ff;
   wire [CONFIG_DW-1:0]                msr_elsa_ff;
   wire [CONFIG_DW*4-1:0]   msr_sr_ff;
   wire                                psr_rm_set;
   wire                                psr_imme_msk;
   wire                                psr_dmme_msk;
   wire                                psr_ire_msk;
   wire                                psr_ld;
   wire                                psr_rm_we;
   wire                                psr_rm_nxt;
   wire                                psr_imme_we;
   wire                                psr_imme_nxt;
   wire                                psr_dmme_we;
   wire                                psr_dmme_nxt;
   wire                                psr_ire_we;
   wire                                psr_ire_nxt;
   wire                                epsr_we;
   wire [10-1:0]             epsr_nxt;
   wire                                epsr_rm_nold;
   wire                                epsr_ire_nold;
   wire                                epsr_imme_nold;
   wire                                epsr_dmme_nold;
   genvar                              i;
   assign psr_ld = msr_psr_save;
   assign psr_rm_set = msr_psr_save;
   assign psr_imme_msk = ~msr_psr_save;
   assign psr_dmme_msk = ~msr_psr_save;
   assign psr_ire_msk = ~msr_psr_save;
   assign epsr_we = (msr_epsr_we | msr_psr_save);
   assign epsr_nxt = msr_psr_save ? msr_psr_nold : msr_epsr_nxt;
   assign psr_rm_we = (msr_psr_rm_we | msr_psr_restore);
   assign psr_rm_nxt = (msr_psr_restore) ? epsr_rm_nold : msr_psr_rm_nxt;
   assign psr_imme_we = (msr_psr_imme_we | msr_psr_restore);
   assign psr_imme_nxt = (msr_psr_restore) ? epsr_imme_nold : msr_psr_imme_nxt;
   assign psr_dmme_we = (msr_psr_dmme_we | msr_psr_restore);
   assign psr_dmme_nxt = (msr_psr_restore) ? epsr_dmme_nold : msr_psr_dmme_nxt;
   assign psr_ire_we = (msr_psr_ire_we | msr_psr_restore);
   assign psr_ire_nxt = (msr_psr_restore) ? epsr_ire_nold : msr_psr_ire_nxt;
   ysyx_20210479_mDFF_lr #(.DW(1), .RST_VECTOR(1'b1)) ff_msr_psr_rm (.CLK(clk), .RST(rst), .LOAD(psr_rm_we|psr_ld), .D(psr_rm_nxt|psr_rm_set), .Q(msr_psr_rm_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_ire (.CLK(clk), .RST(rst), .LOAD(psr_ire_we|psr_ld), .D(psr_ire_nxt&psr_ire_msk), .Q(msr_psr_ire_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_imme (.CLK(clk), .RST(rst), .LOAD(psr_imme_we|psr_ld), .D(psr_imme_nxt&psr_imme_msk), .Q(msr_psr_imme_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_dmme (.CLK(clk), .RST(rst), .LOAD(psr_dmme_we|psr_ld), .D(psr_dmme_nxt&psr_dmme_msk), .Q(msr_psr_dmme_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_ice (.CLK(clk), .RST(rst), .LOAD(msr_psr_ice_we), .D(msr_psr_ice_nxt), .Q(msr_psr_ice_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_dce (.CLK(clk), .RST(rst), .LOAD(msr_psr_dce_we), .D(msr_psr_dce_nxt), .Q(msr_psr_dce_ff) );
   ysyx_20210479_mDFF_lr #(.DW(10)) ff_msr_epsr (.CLK(clk), .RST(rst), .LOAD(epsr_we), .D(epsr_nxt), .Q(msr_epsr_ff) );
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_DW)) ff_msr_epc (.CLK(clk), .RST(rst), .LOAD(msr_epc_we), .D(msr_epc_nxt), .Q(msr_epc_ff) );
   ysyx_20210479_mDFF_lr #(.DW(CONFIG_DW)) dff_msr_elsa (.CLK(clk), .RST(rst), .LOAD(msr_elsa_we), .D(msr_elsa_nxt), .Q(msr_elsa_ff) );
   generate
      for(i=0;i<4;i=i+1)
         ysyx_20210479_mDFF_l #(.DW(CONFIG_DW)) dff_sr (.CLK(clk), .LOAD(msr_sr_we[i]), .D(msr_sr_nxt), .Q(msr_sr_ff[i*CONFIG_DW +: CONFIG_DW]) );
   endgenerate
   assign msr_psr_rm = (psr_rm_we|psr_ld) ? (psr_rm_nxt|psr_rm_set) : msr_psr_rm_ff;
   assign msr_psr_ire = (psr_ire_we|psr_ld) ? (psr_ire_nxt&psr_ire_msk) : msr_psr_ire_ff;
   assign msr_psr_imme = (psr_imme_we|psr_ld) ? (psr_imme_nxt&psr_imme_msk) : msr_psr_imme_ff;
   assign msr_psr_dmme = (psr_dmme_we|psr_ld) ? (psr_dmme_nxt&psr_dmme_msk) : msr_psr_dmme_ff;
   assign msr_psr_rm_nold = (psr_rm_we) ? psr_rm_nxt : msr_psr_rm_ff;
   assign msr_psr_ire_nold = (psr_ire_we) ? psr_ire_nxt : msr_psr_ire_ff;
   assign msr_psr_imme_nold = (psr_imme_we) ? psr_imme_nxt : msr_psr_imme_ff;
   assign msr_psr_dmme_nold = (psr_dmme_we) ? psr_dmme_nxt : msr_psr_dmme_ff;
   assign msr_psr_ice = (msr_psr_ice_we) ? (msr_psr_ice_nxt) : msr_psr_ice_ff;
   assign msr_psr_dce = (msr_psr_dce_we) ? (msr_psr_dce_nxt) : msr_psr_dce_ff;
   assign msr_epsr = epsr_we ? epsr_nxt : msr_epsr_ff;
   assign msr_epc = msr_epc_we ? msr_epc_nxt : msr_epc_ff;
   assign msr_elsa = msr_elsa_we ? msr_elsa_nxt : msr_elsa_ff;
   generate
      for(i=0;i<4;i=i+1)
         assign msr_sr[i*CONFIG_DW +: CONFIG_DW] = (msr_sr_we[i]) ? msr_sr_nxt : msr_sr_ff[i*CONFIG_DW +: CONFIG_DW];
   endgenerate
   assign msr_psr = {msr_psr_dce,msr_psr_ice,msr_psr_dmme,msr_psr_imme,msr_psr_ire,msr_psr_rm,1'b0,1'b0,1'b0,1'b0};
   assign msr_psr_nold = {msr_psr_dce,msr_psr_ice,msr_psr_dmme_nold,msr_psr_imme_nold,msr_psr_ire_nold,msr_psr_rm_nold,1'b0,1'b0,1'b0,1'b0};
   assign {epsr_dmme_nold,epsr_imme_nold,epsr_ire_nold,epsr_rm_nold} = msr_epsr_ff[7:4];
   assign msr_cpuid = {{CONFIG_DW-26{1'b0}},CPUID_FTSC,CPUID_FIRQC,CPUID_FFPU,CPUID_FDBG,CPUID_FDCA,CPUID_FICA,CPUID_FDMM,CPUID_FIMM,CPUID_REV[9:0],CPUID_VER[7:0]};
   assign msr_coreid = {CONFIG_DW{1'b0}};
endmodule
module ysyx_20210479_frontend
#(
   parameter                           CONFIG_AW = 32,
   parameter                           CONFIG_DW = 32,
   parameter                           CONFIG_P_FETCH_WIDTH = 1,
   parameter                           CONFIG_P_ISSUE_WIDTH = 1,
   parameter                           CONFIG_P_IQ_DEPTH = 4,
   parameter                           CONFIG_P_PAGE_SIZE = 13,
   parameter                           CONFIG_ITLB_P_SETS = 0,
   parameter                           CONFIG_IC_P_LINE = 6,
   parameter                           CONFIG_IC_P_SETS = 6,
   parameter                           CONFIG_IC_P_WAYS = 2,
   parameter                           CONFIG_PHT_P_NUM = 9,
   parameter                           CONFIG_BTB_P_NUM = 9,
   parameter [CONFIG_AW-1:0]           CONFIG_ERST_VECTOR = 0,
   parameter                           CONFIG_IMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           AXI_P_DW_BYTES = 3,
   parameter                           AXI_UNCACHED_P_DW_BYTES = 2,
   parameter                           AXI_ADDR_WIDTH = 64,
   parameter                           AXI_ID_WIDTH = 4,
   parameter                           AXI_USER_WIDTH = 1
)
(
   input                               clk,
   input                               rst,
   input                               flush,
   input [(CONFIG_AW-2 )-1:0]                   flush_tgt,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_valid,
   input [CONFIG_P_ISSUE_WIDTH:0]      id_pop_cnt,
   output [((2 <<1)*8) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_ins,
   output [(CONFIG_AW-2 ) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_pc,
   output [2 * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_exc,
   output [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_bpu_upd,
   input                               bpu_wb,
   input                               bpu_wb_is_bcc,
   input                               bpu_wb_is_breg,
   input                               bpu_wb_is_brel,
   input                               bpu_wb_taken,
   input [(CONFIG_AW-2 )-1:0]                   bpu_wb_pc,
   input [(CONFIG_AW-2 )-1:0]                   bpu_wb_npc_act,
   input [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]              bpu_wb_upd,
   input                               msr_psr_imme,
   input                               msr_psr_rm,
   input                               msr_psr_ice,
   output [CONFIG_DW-1:0]              msr_immid,
   input [CONFIG_ITLB_P_SETS-1:0]      msr_imm_tlbl_idx,
   input [CONFIG_DW-1:0]               msr_imm_tlbl_nxt,
   input                               msr_imm_tlbl_we,
   input [CONFIG_ITLB_P_SETS-1:0]      msr_imm_tlbh_idx,
   input [CONFIG_DW-1:0]               msr_imm_tlbh_nxt,
   input                               msr_imm_tlbh_we,
   output [CONFIG_DW-1:0]              msr_icid,
   input [CONFIG_DW-1:0]               msr_icinv_nxt,
   input                               msr_icinv_we,
   output                              msr_icinv_ready,
   input                               ibus_ARREADY,
   output                              ibus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         ibus_ARADDR,
   output [2:0]                        ibus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           ibus_ARID,
   output [AXI_USER_WIDTH-1:0]         ibus_ARUSER,
   output [7:0]                        ibus_ARLEN,
   output [2:0]                        ibus_ARSIZE,
   output [1:0]                        ibus_ARBURST,
   output                              ibus_ARLOCK,
   output [3:0]                        ibus_ARCACHE,
   output [3:0]                        ibus_ARQOS,
   output [3:0]                        ibus_ARREGION,
   output                              ibus_RREADY,
   input                               ibus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  ibus_RDATA,
   input  [1:0]                        ibus_RRESP,
   input                               ibus_RLAST,
   input  [AXI_ID_WIDTH-1:0]           ibus_RID,
   input  [AXI_USER_WIDTH-1:0]         ibus_RUSER
);
   localparam P_FETCH_DW_BYTES         = (2  + CONFIG_P_FETCH_WIDTH);
   localparam FW                       = (1<<CONFIG_P_FETCH_WIDTH);
   wire                 ic_stall_req;           
   wire [((2 <<1)*8)*(1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_ins;
   wire                 iq_ready;               
   wire                                p_ce;
   wire [CONFIG_P_PAGE_SIZE-1:0]       vpo;
   wire                                pred_branch_taken;
   wire [(CONFIG_AW-2 )-1:0]                    pred_branch_tgt;
   wire [CONFIG_AW-1:0]                pc;
   reg [CONFIG_AW-1:0]                 pc_nxt;
   wire [CONFIG_AW-1:0]                s1i_fetch_vaddr;
   wire [FW-1:0]                       s1i_fetch_aligned;
   wire [(CONFIG_AW-2 )-1:0]                    s1i_pc                           [FW-1:0];
   wire [(CONFIG_AW-2 )*FW-1:0]                 s1i_bpu_pc;
   wire [CONFIG_P_FETCH_WIDTH:0]       s1i_push_offset;
   wire [(CONFIG_AW-2 )-1:0]                    s1o_pc                           [FW-1:0];
   wire [2-1:0]               s1o_exc;
   wire [FW-1:0]                       s1o_fetch_aligned;
   wire [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] s1o_tlb_ppn;
   wire                                s1o_tlb_uncached;
   wire                                s1o_msr_psr_ice;
   wire                                s2i_kill_req;
   wire                                s2i_uncached;
   wire [CONFIG_P_FETCH_WIDTH:0]       s1o_push_cnt;
   wire [CONFIG_P_FETCH_WIDTH:0]       s1o_push_offset;
   wire [(CONFIG_AW-2 )*FW-1:0]                 s1o_bpu_npc_packed;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*FW-1:0]            s1o_bpu_upd_packed;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]               s1o_bpu_upd                      [FW-1:0];
   wire [FW-1:0]                       s1o_bpu_taken;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]               s2i_bpu_upd                      [FW-1:0];
   reg [FW-1:0]                        s2i_valid_msk;
   wire [(CONFIG_AW-2 )-1:0]                    s2o_pc                           [FW-1:0];
   wire [2-1:0]               s2o_exc;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]               s2o_bpu_upd                      [FW-1:0];
   wire                                s2o_valid;
   wire [CONFIG_P_FETCH_WIDTH:0]       s2o_push_cnt;
   wire [CONFIG_P_FETCH_WIDTH:0]       s2o_push_offset;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_bpu_upd;
   wire [2*(1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_exc;
   wire [(CONFIG_AW-2 )*(1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_pc;
   wire [CONFIG_P_FETCH_WIDTH:0] iq_push_cnt;  
   wire [CONFIG_P_FETCH_WIDTH:0] iq_push_offset;
   genvar i;
   integer j;
   ysyx_20210479_icache
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_IC_P_LINE               (CONFIG_IC_P_LINE),
        .CONFIG_IC_P_SETS               (CONFIG_IC_P_SETS),
        .CONFIG_IC_P_WAYS               (CONFIG_IC_P_WAYS),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_UNCACHED_P_DW_BYTES        (AXI_UNCACHED_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_I_CACHE
      (
       .stall_req                       (ic_stall_req),          
       .ins                             (iq_ins[((2 <<1)*8)*(1<<CONFIG_P_FETCH_WIDTH)-1:0]), 
       .valid                           (s2o_valid),             
       .msr_icid                        (msr_icid[CONFIG_DW-1:0]),
       .msr_icinv_ready                 (msr_icinv_ready),
       .ibus_ARVALID                    (ibus_ARVALID),
       .ibus_ARADDR                     (ibus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .ibus_ARPROT                     (ibus_ARPROT[2:0]),
       .ibus_ARID                       (ibus_ARID[AXI_ID_WIDTH-1:0]),
       .ibus_ARUSER                     (ibus_ARUSER[AXI_USER_WIDTH-1:0]),
       .ibus_ARLEN                      (ibus_ARLEN[7:0]),
       .ibus_ARSIZE                     (ibus_ARSIZE[2:0]),
       .ibus_ARBURST                    (ibus_ARBURST[1:0]),
       .ibus_ARLOCK                     (ibus_ARLOCK),
       .ibus_ARCACHE                    (ibus_ARCACHE[3:0]),
       .ibus_ARQOS                      (ibus_ARQOS[3:0]),
       .ibus_ARREGION                   (ibus_ARREGION[3:0]),
       .ibus_RREADY                     (ibus_RREADY),
       .clk                             (clk),
       .rst                             (rst),
       .vpo                             (vpo[CONFIG_P_PAGE_SIZE-1:0]),
       .ppn_s2                          (s1o_tlb_ppn),           
       .uncached_s2                     (s2i_uncached),          
       .kill_req_s2                     (s2i_kill_req),          
       .msr_icinv_nxt                   (msr_icinv_nxt[CONFIG_DW-1:0]),
       .msr_icinv_we                    (msr_icinv_we),
       .ibus_ARREADY                    (ibus_ARREADY),
       .ibus_RVALID                     (ibus_RVALID),
       .ibus_RDATA                      (ibus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .ibus_RLAST                      (ibus_RLAST),
       .ibus_RRESP                      (ibus_RRESP[1:0]),
       .ibus_RID                        (ibus_RID[AXI_ID_WIDTH-1:0]),
       .ibus_RUSER                      (ibus_RUSER[AXI_USER_WIDTH-1:0]));
   ysyx_20210479_bpu
      #(
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH))
   U_BPU
      (
         .clk                           (clk),
         .rst                           (rst),
         .re                            (p_ce),
         .valid                         (s1o_fetch_aligned),
         .pc                            (s1i_bpu_pc),
         .npc                           (s1o_bpu_npc_packed),
         .upd                           (s1o_bpu_upd_packed),
         .bpu_wb                        (bpu_wb),
         .bpu_wb_is_bcc                 (bpu_wb_is_bcc),
         .bpu_wb_is_breg                (bpu_wb_is_breg),
         .bpu_wb_is_brel                (bpu_wb_is_brel),
         .bpu_wb_taken                  (bpu_wb_taken),
         .bpu_wb_pc                     (bpu_wb_pc),
         .bpu_wb_npc_act                (bpu_wb_npc_act),
         .bpu_wb_upd                    (bpu_wb_upd)
      );
   ysyx_20210479_immu
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_IMMU_ENABLE_UNCACHED_SEG(CONFIG_IMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_ITLB_P_SETS             (CONFIG_ITLB_P_SETS))
   U_I_MMU
      (
         .clk                             (clk),
         .rst                             (rst),
         .re                              (p_ce),
         .vpn                             (s1i_fetch_vaddr[CONFIG_P_PAGE_SIZE +: CONFIG_AW-CONFIG_P_PAGE_SIZE]),
         .ppn                             (s1o_tlb_ppn),
         .EITM                            (s1o_exc[0]),
         .EIPF                            (s1o_exc[1]),
         .uncached                        (s1o_tlb_uncached),
         .msr_psr_imme                    (msr_psr_imme),
         .msr_psr_rm                      (msr_psr_rm),
         .msr_immid                       (msr_immid),
         .msr_imm_tlbl_idx                (msr_imm_tlbl_idx),
         .msr_imm_tlbl_nxt                (msr_imm_tlbl_nxt),
         .msr_imm_tlbl_we                 (msr_imm_tlbl_we),
         .msr_imm_tlbh_idx                (msr_imm_tlbh_idx),
         .msr_imm_tlbh_nxt                (msr_imm_tlbh_nxt),
         .msr_imm_tlbh_we                 (msr_imm_tlbh_we)
      );
   assign s2i_kill_req = (|s1o_exc);
   assign s2i_uncached = (s1o_tlb_uncached | ~s1o_msr_psr_ice);
   generate
      for(i=0;i<FW;i=i+1)
         begin
            assign s1i_bpu_pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )] = s1i_pc[i];
            assign s1o_bpu_upd[i] = s1o_bpu_upd_packed[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)];
            assign s1o_bpu_taken[i] = s1o_bpu_upd[i][0];
         end
   endgenerate
   always @(*)
      begin
         s2i_valid_msk[0] = 'b1;
         for(j=1;j<FW;j=j+1)
            s2i_valid_msk[j] = s2i_valid_msk[j-1] & ~s1o_bpu_taken[j-1];
      end
   generate
      for(i=0;i<FW;i=i+1)
         assign s1i_fetch_aligned[i] = (pc_nxt[2  +: CONFIG_P_FETCH_WIDTH] <= i);
   endgenerate
   ysyx_20210479_pmux_v #(.SELW(FW), .DW((CONFIG_AW-2 ))) pmux_s1o_bpu_npc (.sel(s1o_bpu_taken), .din(s1o_bpu_npc_packed), .dout(pred_branch_tgt), .valid(pred_branch_taken) );
   always @(*)
      if (flush)
         pc_nxt = {flush_tgt, {2 {1'b0}}};
      else if (~p_ce)
         pc_nxt = pc;
      else if (pred_branch_taken)
         pc_nxt = {pred_branch_tgt, {2 {1'b0}}};
      else
         pc_nxt = pc + {{CONFIG_AW-CONFIG_P_FETCH_WIDTH-1-2 {1'b0}}, s1o_push_cnt, {2 {1'b0}}};
   ysyx_20210479_mDFF_r # (.DW(CONFIG_AW), .RST_VECTOR(CONFIG_ERST_VECTOR)) ff_pc (.CLK(clk), .RST(rst), .D(pc_nxt), .Q(pc) );
   assign p_ce = (~ic_stall_req & iq_ready);
   assign s1i_fetch_vaddr = {pc_nxt[CONFIG_AW-1:P_FETCH_DW_BYTES], {P_FETCH_DW_BYTES{1'b0}}}; 
   ysyx_20210479_popcnt #(.DW(FW), .P_DW(CONFIG_P_FETCH_WIDTH)) popc_1 (.bitmap(~s1i_fetch_aligned), .count(s1i_push_offset) );
   ysyx_20210479_popcnt #(.DW(FW), .P_DW(CONFIG_P_FETCH_WIDTH)) popc_2 (.bitmap(s1o_fetch_aligned & s2i_valid_msk), .count(s1o_push_cnt) );
   assign vpo = s1i_fetch_vaddr[CONFIG_P_PAGE_SIZE-1:0];
   ysyx_20210479_mDFF_lr # (.DW(FW)) ff_s1o_fetch_aligned (.CLK(clk), .RST(rst), .LOAD(p_ce|flush), .D(s1i_fetch_aligned & {FW{~flush}}), .Q(s1o_fetch_aligned) );
   ysyx_20210479_mDFF_lr # (.DW(CONFIG_P_FETCH_WIDTH+1)) ff_s2o_push_cnt (.CLK(clk), .RST(rst), .LOAD(p_ce|flush), .D(s1o_push_cnt & {CONFIG_P_FETCH_WIDTH+1{~flush}}), .Q(s2o_push_cnt) );
   ysyx_20210479_mDFF_lr # (.DW(2)) ff_s2o_exc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_exc), .Q(s2o_exc) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_msr_psr_ice (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(msr_psr_ice), .Q(s1o_msr_psr_ice) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_P_FETCH_WIDTH+1)) ff_s1o_push_offset (.CLK(clk), .LOAD(p_ce), .D(s1i_push_offset), .Q(s1o_push_offset) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_P_FETCH_WIDTH+1)) ff_s2o_push_offset (.CLK(clk), .LOAD(p_ce), .D(s1o_push_offset), .Q(s2o_push_offset) );
   generate
      for(i=0;i<FW;i=i+1)
         begin
            assign s1i_pc[i] = (pc_nxt[CONFIG_AW-1: 2 ] + i - {{(CONFIG_AW-2 )-CONFIG_P_FETCH_WIDTH-1{1'b0}}, s1i_push_offset});
            ysyx_20210479_mDFF_lr # (.DW((CONFIG_AW-2 ))) ff_s1o_pc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1i_pc[i]), .Q(s1o_pc[i]) );
            ysyx_20210479_mDFF_lr # (.DW((CONFIG_AW-2 ))) ff_s2o_pc (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_pc[i]), .Q(s2o_pc[i]) );
            ysyx_20210479_mDFF_lr # (.DW((2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1))) ff_s2o_bpu_upd (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_bpu_upd[i]), .Q(s2o_bpu_upd[i]) );
            assign iq_pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )] = s2o_pc[i];
            assign iq_exc[i*2 +: 2] = s2o_exc;
            assign iq_bpu_upd[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)] = s2o_bpu_upd[i];
         end
   endgenerate
   assign iq_push_cnt = (s2o_push_cnt & {CONFIG_P_FETCH_WIDTH+1{s2o_valid & p_ce}});
   assign iq_push_offset = (s2o_push_offset);
   ysyx_20210479_prefetch_buf
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH),
        .CONFIG_P_IQ_DEPTH              (CONFIG_P_IQ_DEPTH),
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM))
   U_PREFETCH_BUF
      (
       .iq_ready                        (iq_ready),
       .id_valid                        (id_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_ins                          (id_ins[((2 <<1)*8)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_pc                           (id_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_exc                          (id_exc[2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_bpu_upd                      (id_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .flush                           (flush),
       .iq_ins                          (iq_ins[((2 <<1)*8)*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
       .iq_pc                           (iq_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
       .iq_exc                          (iq_exc[2*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
       .iq_bpu_upd                      (iq_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_FETCH_WIDTH)-1:0]),
       .iq_push_cnt                     (iq_push_cnt[CONFIG_P_FETCH_WIDTH:0]),
       .iq_push_offset                  (iq_push_offset[CONFIG_P_FETCH_WIDTH:0]),
       .id_pop_cnt                      (id_pop_cnt[CONFIG_P_ISSUE_WIDTH:0]));
endmodule
module ysyx_20210479_icache
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_FETCH_WIDTH = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_IC_P_LINE = 0,
   parameter                           CONFIG_IC_P_SETS = 0,
   parameter                           CONFIG_IC_P_WAYS = 0,
   parameter                           AXI_P_DW_BYTES  = 3,
   parameter                           AXI_UNCACHED_P_DW_BYTES = 2,
   parameter                           AXI_ADDR_WIDTH    = 64,
   parameter                           AXI_ID_WIDTH      = 4,
   parameter                           AXI_USER_WIDTH    = 1
)
(
   input                               clk,
   input                               rst,
   output                              stall_req,
   input [CONFIG_P_PAGE_SIZE-1:0]      vpo,
   input [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] ppn_s2,
   input                               uncached_s2,
   input                               kill_req_s2,
   output [((2 <<1)*8) * (1<<CONFIG_P_FETCH_WIDTH)-1:0] ins,
   output                              valid,
   output [CONFIG_DW-1:0]              msr_icid,
   input [CONFIG_DW-1:0]               msr_icinv_nxt,
   input                               msr_icinv_we,
   output                              msr_icinv_ready,
   input                               ibus_ARREADY,
   output                              ibus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         ibus_ARADDR,
   output [2:0]                        ibus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           ibus_ARID,
   output [AXI_USER_WIDTH-1:0]         ibus_ARUSER,
   output [7:0]                        ibus_ARLEN,
   output [2:0]                        ibus_ARSIZE,
   output [1:0]                        ibus_ARBURST,
   output                              ibus_ARLOCK,
   output [3:0]                        ibus_ARCACHE,
   output [3:0]                        ibus_ARQOS,
   output [3:0]                        ibus_ARREGION,
   output                              ibus_RREADY,
   input                               ibus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  ibus_RDATA,
   input                               ibus_RLAST,
   input  [1:0]                        ibus_RRESP, 
   input  [AXI_ID_WIDTH-1:0]           ibus_RID, 
   input  [AXI_USER_WIDTH-1:0]         ibus_RUSER 
);
   localparam TAG_WIDTH                = (CONFIG_AW - CONFIG_IC_P_SETS - CONFIG_IC_P_LINE);
   localparam TAG_V_RAM_AW             = (CONFIG_IC_P_SETS);
   localparam TAG_V_RAM_DW             = (TAG_WIDTH + 1); 
   localparam PAYLOAD_DW               = (((2 <<1)*8) * (1<<CONFIG_P_FETCH_WIDTH));
   localparam PAYLOAD_P_DW_BYTES       = (2  + CONFIG_P_FETCH_WIDTH); 
   localparam PAYLOAD_AW               = (CONFIG_IC_P_SETS + CONFIG_IC_P_LINE - PAYLOAD_P_DW_BYTES);
   localparam AXI_FETCH_SIZE           = (PAYLOAD_P_DW_BYTES <= AXI_P_DW_BYTES) ? PAYLOAD_P_DW_BYTES : AXI_P_DW_BYTES;
   localparam AXI_UNCACHED_DW          = (1<<AXI_UNCACHED_P_DW_BYTES)*8;
   reg [CONFIG_IC_P_SETS-1:0]          s1i_line_addr;
   reg [TAG_V_RAM_DW-1:0]              s1i_replace_tag_v;
   wire                                s1i_tag_v_re;
   wire                                s1i_tag_v_we            [(1<<CONFIG_IC_P_WAYS)-1:0];
   wire                                s1i_payload_re;
   reg [PAYLOAD_AW-1:0]                s1i_payload_addr;
   wire [PAYLOAD_DW/8-1:0]             s1i_payload_we          [(1<<CONFIG_IC_P_WAYS)-1:0];
   wire [PAYLOAD_DW-1:0]               s1i_payload_din;
   wire [AXI_UNCACHED_DW/8-1:0]        s1i_uncached_align_we;
   wire [AXI_UNCACHED_DW-1:0]          s1i_uncached_align_din;
   wire [PAYLOAD_DW/8-1:0]             s1i_uncached_we;
   wire [PAYLOAD_DW-1:0]               s1i_uncached_din;
   wire [PAYLOAD_DW/8-1:0]             s1i_payload_tgt_we;
   wire [CONFIG_IC_P_SETS-1:0]         s1o_line_addr;
   wire [PAYLOAD_AW-1:0]               s1o_payload_addr;
   wire                                s1o_valid;
   wire [PAYLOAD_DW*(1<<CONFIG_IC_P_WAYS)-1:0] s1o_payload;
   wire [PAYLOAD_DW-1:0]               s1o_match_payload;
   wire [TAG_V_RAM_DW-1:0]             s1o_tag_v               [(1<<CONFIG_IC_P_WAYS)-1:0];
   wire [CONFIG_P_PAGE_SIZE-1:0]       s1o_vpo;
   wire [CONFIG_AW-1:0]                s2i_paddr;
   wire [TAG_WIDTH-1:0]                s2i_tag                 [(1<<CONFIG_IC_P_WAYS)-1:0];
   wire                                s2i_v                   [(1<<CONFIG_IC_P_WAYS)-1:0];
   wire [(1<<CONFIG_IC_P_WAYS)-1:0]    s2i_hit_vec;
   wire                                s2i_hit;
   wire                                s2i_refill_get_dat;
   wire                                s2i_uncached_get_dat;
   reg [PAYLOAD_DW-1:0]                s2i_ins;
   wire [CONFIG_AW-1:0]                s1o_op_inv_paddr;
   wire [CONFIG_IC_P_SETS-1:0]         s2o_line_addr;
   wire                                s2o_valid;
   wire [CONFIG_AW-1:0]                s2o_paddr;
   wire [(1<<CONFIG_IC_P_WAYS)-1:0]    s2o_fsm_free_way;
   reg [2:0]                           fsm_state_nxt;
   wire [2:0]                          fsm_state_ff;
   wire [(1<<CONFIG_IC_P_WAYS)-1:0]    fsm_free_way, fsm_free_way_nxt;
   wire [CONFIG_IC_P_SETS-1:0]         fsm_boot_cnt;
   wire [CONFIG_IC_P_SETS:0]           fsm_boot_cnt_nxt_carry;
   wire [CONFIG_IC_P_LINE-1:0]         fsm_refill_cnt;
   reg [CONFIG_IC_P_LINE-1:0]          fsm_refill_cnt_nxt;
   wire [PAYLOAD_P_DW_BYTES-1:0]       fsm_uncached_cnt;
   reg [PAYLOAD_P_DW_BYTES-1:0]        fsm_uncached_cnt_nxt;
   wire [PAYLOAD_P_DW_BYTES:0]         fsm_uncached_cnt_nxt_carry;
   reg                                 fsm_uncached_rd_req;
   wire                                p_ce;
   wire                                ar_set, ar_clr;
   wire                                hds_axi_R;
   wire                                hds_axi_R_last;
   wire [CONFIG_AW-1:0]                axi_paddr_nxt;
   wire [AXI_ADDR_WIDTH-1:0]           axi_ar_addr_nxt;
   localparam [2:0] S_BOOT             = 3'd0;
   localparam [2:0] S_IDLE             = 3'd1;
   localparam [2:0] S_REPLACE          = 3'd2;
   localparam [2:0] S_REFILL           = 3'd3;
   localparam [2:0] S_INVALIDATE       = 3'd4;
   localparam [2:0] S_RELOAD_S1O       = 3'd5;
   localparam [2:0] S_UNCACHED_BOOT    = 3'd6;
   localparam [2:0] S_UNCACHED_READ    = 3'd7;
   genvar way, i, j;
   assign p_ce = (~stall_req);
   assign s2i_paddr = {ppn_s2, s1o_vpo};
   generate
      for(way=0; way<(1<<CONFIG_IC_P_WAYS); way=way+1)
         begin : gen_ways
            ysyx_20210479_mRAM_s_s_be
               #(
                  .P_DW (PAYLOAD_P_DW_BYTES + 3),
                  .AW   (PAYLOAD_AW)
               )
            U_PAYLOAD_RAM
               (
                  .CLK  (clk),
                  .ADDR (s1i_payload_addr),
                  .RE   (s1i_payload_re),
                  .DOUT (s1o_payload[way*PAYLOAD_DW +: PAYLOAD_DW]),
                  .WE   (s1i_payload_we[way]),
                  .DIN  (s1i_payload_din)
               );
            ysyx_20210479_mRF_1wr
               #(
                  .DW   (TAG_V_RAM_DW),
                  .AW   (TAG_V_RAM_AW)
               )
            U_TAG_V_RAM
               (
                  .CLK  (clk),
                  .ADDR (s1i_line_addr),
                  .RE   (s1i_tag_v_re),
                  .RDATA (s1o_tag_v[way]),
                  .WE   (s1i_tag_v_we[way]),
                  .WDATA (s1i_replace_tag_v)
               );
            assign {s2i_tag[way], s2i_v[way]} = s1o_tag_v[way];
            assign s2i_hit_vec[way] = (s2i_v[way] & (s2i_tag[way] == s2i_paddr[CONFIG_AW-1:CONFIG_IC_P_LINE+CONFIG_IC_P_SETS]) );
         end
   endgenerate
   ysyx_20210479_pmux_v #(.SELW(1<<CONFIG_IC_P_WAYS), .DW(PAYLOAD_DW)) pmux_s1o_payload (.sel(s2i_hit_vec), .din(s1o_payload), .dout(s1o_match_payload), .valid(s2i_hit) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s1o_valid (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(1'b1), .Q(s1o_valid) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_P_PAGE_SIZE)) ff_s1o_vpo (.CLK(clk), .LOAD(p_ce), .D(vpo), .Q(s1o_vpo) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_AW)) ff_s1o_op_inv_paddr (.CLK(clk), .LOAD(p_ce), .D(msr_icinv_nxt), .Q(s1o_op_inv_paddr) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_IC_P_SETS)) ff_s1o_line_addr (.CLK(clk), .LOAD(p_ce), .D(s1i_line_addr), .Q(s1o_line_addr) );
   ysyx_20210479_mDFF_l # (.DW(PAYLOAD_AW)) ff_s1o_payload_addr (.CLK(clk), .LOAD(p_ce), .D(s1i_payload_addr), .Q(s1o_payload_addr) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_IC_P_SETS)) ff_s2o_line_addr (.CLK(clk), .LOAD(p_ce), .D(s1o_line_addr), .Q(s2o_line_addr) );
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_s2o_valid (.CLK(clk), .RST(rst), .LOAD(p_ce), .D(s1o_valid), .Q(s2o_valid) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_AW)) ff_s2o_paddr (.CLK(clk), .LOAD(p_ce), .D(s2i_paddr), .Q(s2o_paddr) );
   always @(*)
      begin
         fsm_state_nxt = fsm_state_ff;
         fsm_uncached_rd_req = 'b0;
         case (fsm_state_ff)
            S_BOOT:
               if (fsm_boot_cnt_nxt_carry[CONFIG_IC_P_SETS])
                  fsm_state_nxt = S_IDLE;
            S_IDLE:
               if (msr_icinv_we) 
                  fsm_state_nxt = S_INVALIDATE;
               else if (s1o_valid & uncached_s2 & ~kill_req_s2) 
                  fsm_state_nxt = S_UNCACHED_BOOT;
               else if (s1o_valid & ~s2i_hit & ~uncached_s2 & ~kill_req_s2) 
                  fsm_state_nxt = S_REPLACE;
            S_REPLACE:
               fsm_state_nxt = S_REFILL;
            S_REFILL:
               if (hds_axi_R_last)
                  fsm_state_nxt = S_RELOAD_S1O;
            S_INVALIDATE:
               fsm_state_nxt = S_IDLE;
            S_RELOAD_S1O:
               fsm_state_nxt = S_IDLE;
            S_UNCACHED_BOOT:
               begin
                  fsm_state_nxt = S_UNCACHED_READ;
                  fsm_uncached_rd_req = 'b1;
               end
            S_UNCACHED_READ:
               if (fsm_uncached_cnt_nxt_carry[PAYLOAD_P_DW_BYTES] & hds_axi_R)
                  fsm_state_nxt = S_IDLE;
               else if (hds_axi_R)
                  fsm_uncached_rd_req = 'b1; 
            default: ;
         endcase
      end
   ysyx_20210479_mDFF_r # (.DW(3), .RST_VECTOR(S_BOOT)) ff_state_r (.CLK(clk), .RST(rst), .D(fsm_state_nxt), .Q(fsm_state_ff) );
   assign fsm_free_way_nxt = (fsm_free_way[(1<<CONFIG_IC_P_WAYS)-1])
                              ? {{(1<<CONFIG_IC_P_WAYS)-1{1'b0}}, 1'b1}
                              : {fsm_free_way[(1<<CONFIG_IC_P_WAYS)-2:0], 1'b0};
   ysyx_20210479_mDFF_r #(.DW(1<<CONFIG_IC_P_WAYS), .RST_VECTOR({{(1<<CONFIG_IC_P_WAYS)-1{1'b0}}, 1'b1}) ) ff_fsm_free_idx
      (.CLK(clk), .RST(rst), .D(fsm_free_way_nxt), .Q(fsm_free_way) );
   assign fsm_boot_cnt_nxt_carry = fsm_boot_cnt + 'b1;
   ysyx_20210479_mDFF_r # (.DW(CONFIG_IC_P_SETS)) ff_fsm_boot_cnt_nxt (.CLK(clk), .RST(rst), .D(fsm_boot_cnt_nxt_carry[CONFIG_IC_P_SETS-1:0]), .Q(fsm_boot_cnt) );
   always @(*)
      if ((fsm_state_ff == S_REFILL) & hds_axi_R)
         fsm_refill_cnt_nxt = fsm_refill_cnt + (1<<AXI_FETCH_SIZE);
      else
         fsm_refill_cnt_nxt = fsm_refill_cnt;
   ysyx_20210479_mDFF_r # (.DW(CONFIG_IC_P_LINE)) ff_fsm_refill_cnt (.CLK(clk), .RST(rst), .D(fsm_refill_cnt_nxt), .Q(fsm_refill_cnt) );
   always @(*)
      if ((fsm_state_ff == S_UNCACHED_READ) & hds_axi_R)
         fsm_uncached_cnt_nxt = fsm_uncached_cnt_nxt_carry[PAYLOAD_P_DW_BYTES-1:0];
      else
         fsm_uncached_cnt_nxt = fsm_uncached_cnt;
   assign fsm_uncached_cnt_nxt_carry = fsm_uncached_cnt + (1<<AXI_UNCACHED_P_DW_BYTES);
   ysyx_20210479_mDFF_r # (.DW(PAYLOAD_P_DW_BYTES)) ff_fsm_uncached_cnt (.CLK(clk), .RST(rst), .D(fsm_uncached_cnt_nxt), .Q(fsm_uncached_cnt) );
   always @(*)
      case (fsm_state_ff)
         S_BOOT:
            s1i_line_addr = fsm_boot_cnt;
         S_INVALIDATE:
            s1i_line_addr = s1o_op_inv_paddr[CONFIG_IC_P_LINE +: CONFIG_IC_P_SETS];
         S_REPLACE:
            s1i_line_addr = s2o_line_addr;
         S_RELOAD_S1O:
            s1i_line_addr = s1o_line_addr;
         default:
            s1i_line_addr = vpo[CONFIG_IC_P_LINE +: CONFIG_IC_P_SETS]; 
      endcase
   always @(*)
      case (fsm_state_ff)
         S_REPLACE:
            s1i_replace_tag_v = {s2o_paddr[CONFIG_AW-1:CONFIG_IC_P_LINE+CONFIG_IC_P_SETS], 1'b1};
         default: 
            s1i_replace_tag_v = 'b0;
      endcase
   assign s1i_tag_v_re = (p_ce | (fsm_state_ff==S_RELOAD_S1O));
   generate
      for(way=0; way<(1<<CONFIG_IC_P_WAYS); way=way+1)
         assign s1i_tag_v_we[way] = (fsm_state_ff==S_BOOT) |
                                    (fsm_state_ff==S_INVALIDATE) |
                                    ((fsm_state_ff==S_REPLACE) & (fsm_free_way[way]));
   endgenerate
   ysyx_20210479_mDFF_l #(.DW(1<<CONFIG_IC_P_WAYS)) ff_s2o_fsm_free_way(.CLK(clk), .LOAD(fsm_state_ff==S_REPLACE), .D(fsm_free_way), .Q(s2o_fsm_free_way));
   always @(*)
      case (fsm_state_ff)
         S_REFILL:
            s1i_payload_addr = {s2o_paddr[CONFIG_IC_P_LINE +: CONFIG_IC_P_SETS], fsm_refill_cnt[PAYLOAD_P_DW_BYTES +: CONFIG_IC_P_LINE-PAYLOAD_P_DW_BYTES]};
         S_RELOAD_S1O:
            s1i_payload_addr = s1o_payload_addr;
         default:
            s1i_payload_addr = vpo[PAYLOAD_P_DW_BYTES +: PAYLOAD_AW]; 
      endcase
   assign s1i_payload_re = s1i_tag_v_re;
   ysyx_20210479_align_r
      #(
         .AXI_P_DW_BYTES               (AXI_P_DW_BYTES),
         .PAYLOAD_P_DW_BYTES           (PAYLOAD_P_DW_BYTES),
         .RAM_AW                       (CONFIG_IC_P_LINE)
      )
   U_ALIGN_R
      (
         .i_axi_RDATA                  (ibus_RDATA),
         .i_ram_we                     (fsm_state_ff == S_REFILL),
         .i_ram_addr                   (fsm_refill_cnt),
         .o_ram_wmsk                   (s1i_payload_tgt_we),
         .o_ram_din                    (s1i_payload_din)
      );
   generate
      for(way=0; way<(1<<CONFIG_IC_P_WAYS); way=way+1)
         assign s1i_payload_we[way] = (s1i_payload_tgt_we & {PAYLOAD_DW/8{s2o_fsm_free_way[way]}});
   endgenerate
   ysyx_20210479_align_r
      #(
         .AXI_P_DW_BYTES               (AXI_P_DW_BYTES),
         .PAYLOAD_P_DW_BYTES           (AXI_UNCACHED_P_DW_BYTES),
         .RAM_AW                       (AXI_ADDR_WIDTH)
      )
   U_ALIGN_R_UNCACHED
      (
         .i_axi_RDATA                  (ibus_RDATA),
         .i_ram_we                     (fsm_state_ff == S_UNCACHED_READ),
         .i_ram_addr                   (ibus_ARADDR),
         .o_ram_wmsk                   (s1i_uncached_align_we),
         .o_ram_din                    (s1i_uncached_align_din)
      );
   generate
      for(j=0;j<PAYLOAD_DW/AXI_UNCACHED_DW;j=j+1)
         begin : gen_align_uncached
            assign s1i_uncached_din[j*AXI_UNCACHED_DW +: AXI_UNCACHED_DW] = s1i_uncached_align_din;
            assign s1i_uncached_we[j*AXI_UNCACHED_DW/8 +: AXI_UNCACHED_DW/8] = s1i_uncached_align_we & {AXI_UNCACHED_DW/8{}};
         end
   endgenerate
   assign stall_req = (fsm_state_ff != S_IDLE);
   assign msr_icinv_ready = (~stall_req); 
   assign s2i_refill_get_dat = (s2o_paddr[PAYLOAD_P_DW_BYTES +: CONFIG_IC_P_LINE-PAYLOAD_P_DW_BYTES] ==
                                 fsm_refill_cnt[PAYLOAD_P_DW_BYTES +: CONFIG_IC_P_LINE-PAYLOAD_P_DW_BYTES]);
   assign s2i_uncached_get_dat = (s2o_paddr[PAYLOAD_P_DW_BYTES +: CONFIG_IC_P_LINE-PAYLOAD_P_DW_BYTES] ==
                                 ibus_ARADDR[PAYLOAD_P_DW_BYTES +: CONFIG_IC_P_LINE-PAYLOAD_P_DW_BYTES]);
   generate
      for(j=0;j<PAYLOAD_DW/8;j=j+1)
         begin : gen_output_inner
            always @(*)
               case (fsm_state_ff)
                  S_REFILL:
                     if (s2i_refill_get_dat & s1i_payload_tgt_we[j])
                        s2i_ins[j*8 +: 8] = s1i_payload_din[j*8 +: 8]; 
                     else
                        s2i_ins[j*8 +: 8] = ins[j*8 +: 8];
                  S_UNCACHED_READ:
                     if (s2i_uncached_get_dat & s1i_uncached_we[j])
                        s2i_ins[j*8 +: 8] = s1i_uncached_din[j*8 +: 8]; 
                     else
                        s2i_ins[j*8 +: 8] = ins[j*8 +: 8];
                  default:
                     s2i_ins[j*8 +: 8] = s1o_match_payload[j*8 +: 8]; 
               endcase
         end
   endgenerate
   ysyx_20210479_mDFF_l # (.DW(PAYLOAD_DW)) ff_ins (.CLK(clk), .LOAD(p_ce|(fsm_state_ff==S_REFILL)|(fsm_state_ff==S_UNCACHED_READ)), .D(s2i_ins), .Q(ins) );
   assign valid = (s2o_valid & ~stall_req);
   assign ibus_ARPROT = 3'b000 | 3'b000 | 3'b000;
   assign ibus_ARID = {AXI_ID_WIDTH{1'b0}};
   assign ibus_ARUSER = {AXI_USER_WIDTH{1'b0}};
   assign ibus_ARLEN = (fsm_state_ff==S_REFILL) ? ((1<<(CONFIG_IC_P_LINE-AXI_FETCH_SIZE))-1) : 'b0;
   assign ibus_ARSIZE = (fsm_state_ff==S_REFILL) ? AXI_FETCH_SIZE : AXI_UNCACHED_P_DW_BYTES;
   assign ibus_ARBURST = 2'b01;
   assign ibus_ARLOCK = 'b0;
   assign ibus_ARCACHE = 4'b0010;
   assign ibus_ARQOS = 'b0;
   assign ibus_ARREGION = 'b0;
   assign ar_set = ((fsm_state_ff==S_REPLACE) | fsm_uncached_rd_req);
   assign ar_clr = (ibus_ARREADY & ibus_ARVALID);
   assign axi_paddr_nxt = (fsm_uncached_rd_req)
                           ? {s2o_paddr[PAYLOAD_P_DW_BYTES +: CONFIG_AW - PAYLOAD_P_DW_BYTES], fsm_uncached_cnt_nxt}
                           : {s2o_paddr[CONFIG_IC_P_LINE +: CONFIG_AW - CONFIG_IC_P_LINE], {CONFIG_IC_P_LINE{1'b0}}};
   generate
      if (AXI_ADDR_WIDTH > CONFIG_AW)
         assign axi_ar_addr_nxt = {{AXI_ADDR_WIDTH-CONFIG_AW{1'b0}}, axi_paddr_nxt};
      else if (AXI_ADDR_WIDTH < CONFIG_AW)
         assign axi_ar_addr_nxt = axi_paddr_nxt[AXI_ADDR_WIDTH-1:0];
      else
         assign axi_ar_addr_nxt = axi_paddr_nxt;
   endgenerate
   ysyx_20210479_mDFF_lr # (.DW(1)) ff_axi_ar_valid (.CLK(clk), .RST(rst), .LOAD(ar_set|ar_clr), .D(ar_set|~ar_clr), .Q(ibus_ARVALID) );
   ysyx_20210479_mDFF_lr # (.DW(AXI_ADDR_WIDTH)) ff_axi_ar_addr (.CLK(clk), .RST(rst), .LOAD(ar_set), .D(axi_ar_addr_nxt), .Q(ibus_ARADDR) );
   assign ibus_RREADY = (fsm_state_ff == S_REFILL) | (fsm_state_ff == S_UNCACHED_READ);
   assign hds_axi_R = (ibus_RVALID & ibus_RREADY);
   assign hds_axi_R_last = (hds_axi_R & ibus_RLAST);
   assign msr_icid[3:0] = CONFIG_IC_P_SETS[3:0];
   assign msr_icid[7:4] = CONFIG_IC_P_LINE[3:0];
   assign msr_icid[11:8] = CONFIG_IC_P_WAYS[3:0];
   assign msr_icid[31:12] = 20'b0;
endmodule
module ysyx_20210479_id
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_ISSUE_WIDTH = 0,
   parameter                           CONFIG_PHT_P_NUM = 0,
   parameter                           CONFIG_BTB_P_NUM = 0,
   parameter                           CONFIG_ENABLE_MUL = 0,
   parameter                           CONFIG_ENABLE_DIV = 0,
   parameter                           CONFIG_ENABLE_DIVU = 0,
   parameter                           CONFIG_ENABLE_MOD = 0,
   parameter                           CONFIG_ENABLE_MODU = 0,
   parameter                           CONFIG_ENABLE_ASR = 0
)
(
   input                               clk,
   input                               rst,
   input                               flush,
   input                               stall,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_valid,
   output [CONFIG_P_ISSUE_WIDTH:0]      id_pop_cnt,
   input [((2 <<1)*8) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_ins,
   input [(CONFIG_AW-2 ) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_pc,
   input [2 * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_exc,
   input [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_bpu_upd,
   input                               irq_async,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0]                ex_valid,
   output [9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_alu_opc_bus,
   output [5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lpu_opc_bus,
   output [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_epu_opc_bus,
   output [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bru_opc_bus,
   output [7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lsu_opc_bus,
   output [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bpu_upd,
   output [(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_pc,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_imm,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand1,
   output [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand2,
   output [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_waddr,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_we,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_wdat,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_we,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_waddr,
   input                               ro_ex_s1_load0,
   input                               ro_ex_s2_load0,
   input                               ro_ex_s3_load0,
   output [(1<<CONFIG_P_ISSUE_WIDTH)*2-1:0] arf_RE,
   output [(1<<CONFIG_P_ISSUE_WIDTH)*2*5-1:0] arf_RADDR,
   input [(1<<CONFIG_P_ISSUE_WIDTH)*2*CONFIG_DW-1:0] arf_RDATA
);
   localparam IW                       = (1<<CONFIG_P_ISSUE_WIDTH);
   wire                                p_ce;
   reg [IW-1:0]                        valid_msk;
   wire [IW-1:0]                       valid;
   wire [IW-1:0]                       single_fu;
   reg [IW-1:0]                        raw_dep;
   wire [9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_alu_opc_bus;
   wire [5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_lpu_opc_bus;
   wire [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_epu_opc_bus;
   wire [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_bru_opc_bus;
   wire [7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_lsu_opc_bus;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] s1i_imm;
   wire [IW-1:0]                       rf_we;
   wire [5*IW-1:0]          rf_waddr;
   wire [IW-1:0]                       rf_rs1_re;
   wire [5-1:0]             rf_rs1_addr                   [IW-1:0];
   wire [IW-1:0]                       rf_rs2_re;
   wire [5-1:0]             rf_rs2_addr                   [IW-1:0];
   wire [IW-1:0]                       s1o_rf_rs2_re;
   wire [CONFIG_DW*2*IW-1:0]           byp_dout;
   wire [CONFIG_DW-1:0]                rop1                          [IW-1:0];
   wire [CONFIG_DW-1:0]                rop2                          [IW-1:0];
   wire [2*IW-1:0]                     raw_dep_load0;
   genvar i;
   integer j, k;
   generate
      for(i=0;i<IW;i=i+1)
         begin : gen_dec
            ysyx_20210479_id_dec
               #(
                 .CONFIG_AW             (CONFIG_AW),
                 .CONFIG_DW             (CONFIG_DW),
                 .CONFIG_ENABLE_MUL     (CONFIG_ENABLE_MUL),
                 .CONFIG_ENABLE_DIV     (CONFIG_ENABLE_DIV),
                 .CONFIG_ENABLE_DIVU    (CONFIG_ENABLE_DIVU),
                 .CONFIG_ENABLE_MOD     (CONFIG_ENABLE_MOD),
                 .CONFIG_ENABLE_MODU    (CONFIG_ENABLE_MODU),
                 .CONFIG_ENABLE_ASR     (CONFIG_ENABLE_ASR))
            U_DEC
               (
                  .id_valid            (id_valid[i]),
                  .id_ins              (id_ins[i*((2 <<1)*8) +: ((2 <<1)*8)]),
                  .id_exc              (id_exc[i*2 +: 2]),
                  .irq_async           (irq_async),
                  .single_fu           (single_fu[i]),
                  .alu_opc_bus         (s1i_alu_opc_bus[i*9  +: 9 ]),
                  .lpu_opc_bus         (s1i_lpu_opc_bus[i*5  +: 5 ]),
                  .epu_opc_bus         (s1i_epu_opc_bus[i*8 +: 8]),
                  .bru_opc_bus         (s1i_bru_opc_bus[i*8 +: 8]),
                  .lsu_opc_bus         (s1i_lsu_opc_bus[i*7 +: 7]),
                  .imm                 (s1i_imm[i*CONFIG_DW +: CONFIG_DW]),
                  .rf_we               (rf_we[i]),
                  .rf_waddr            (rf_waddr[i*5 +:5 ]),
                  .rf_rs1_re           (rf_rs1_re[i]),
                  .rf_rs1_addr         (rf_rs1_addr[i]),
                  .rf_rs2_re           (rf_rs2_re[i]),
                  .rf_rs2_addr         (rf_rs2_addr[i])
               );
         end
   endgenerate
   always @(*)
      for(k=0;k<IW;k=k+1)
         begin
            raw_dep[k] = (raw_dep_load0[(k<<1)] | raw_dep_load0[(k<<1)+1]);
            for(j=0;j<k;j=j+1)
               raw_dep[k] = raw_dep[k] | (rf_we[j] &
                                          ((rf_rs1_re[k] & (rf_rs1_addr[k]==rf_waddr[j*5 +:5 ])) |
                                             (rf_rs2_re[k] & (rf_rs2_addr[k]==rf_waddr[j*5 +:5 ]))));
         end
   always @(*)
      begin
         valid_msk[0] = ~raw_dep[0];
         for(j=1;j<IW;j=j+1)
            valid_msk[j] = valid_msk[j-1] & ~single_fu[j] & ~raw_dep[j];
      end
   assign valid = (valid_msk & id_valid);
   ysyx_20210479_popcnt #(.DW(IW), .P_DW(CONFIG_P_ISSUE_WIDTH)) U_CLO (.bitmap(valid & {IW{p_ce}}), .count(id_pop_cnt) );
   assign p_ce = (~stall);
   ysyx_20210479_id_ro
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH))
   U_RO
      (
       .byp_dout                        (byp_dout[CONFIG_DW*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .raw_dep_load0                   (raw_dep_load0[2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .clk                             (clk),
       .ro_ex_s1_rf_dout                (ro_ex_s1_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_dout                (ro_ex_s2_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_dout                (ro_ex_s3_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_wdat                  (ro_cmt_rf_wdat[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_we                  (ro_ex_s1_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_we                  (ro_ex_s2_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_we                  (ro_ex_s3_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_we                    (ro_cmt_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_waddr               (ro_ex_s1_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_waddr               (ro_ex_s2_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_waddr               (ro_ex_s3_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_waddr                 (ro_cmt_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_load0                  (ro_ex_s1_load0),
       .ro_ex_s2_load0                  (ro_ex_s2_load0),
       .ro_ex_s3_load0                  (ro_ex_s3_load0),
       .raddr                           (arf_RADDR[5*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]), 
       .re                              (arf_RE[2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]), 
       .rf_din                          (arf_RDATA[CONFIG_DW*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0])); 
   generate
      for(i=0;i<IW;i=i+1)
         begin
            assign arf_RE[(i<<1)] = (p_ce & rf_rs1_re[i]);
            assign arf_RE[(i<<1)+1] = (p_ce & rf_rs2_re[i]);
            assign arf_RADDR[(i<<1)*5 +: 5] = rf_rs1_addr[i];
            assign arf_RADDR[((i<<1)+1)*5 +: 5] = rf_rs2_addr[i];
            assign rop1[i] = byp_dout[(i<<1)*CONFIG_DW +: CONFIG_DW];
            assign rop2[i] = byp_dout[((i<<1)+1)*CONFIG_DW +: CONFIG_DW];
            assign ex_operand1[i*CONFIG_DW +: CONFIG_DW] = rop1[i];
            assign ex_operand2[i*CONFIG_DW +: CONFIG_DW] = (s1o_rf_rs2_re[i]) ? rop2[i] : ex_imm[i*CONFIG_DW +: CONFIG_DW];
         end
   endgenerate
   ysyx_20210479_mDFF_lr # (.DW(IW)) ff_ex_valid (.CLK(clk), .RST(rst), .LOAD(p_ce|flush), .D(valid & {IW{~flush}}), .Q(ex_valid) );
   ysyx_20210479_mDFF_l # (.DW(9 *IW)) ff_ex_alu_opc_bus (.CLK(clk), .LOAD(p_ce), .D(s1i_alu_opc_bus), .Q(ex_alu_opc_bus) );
   ysyx_20210479_mDFF_l # (.DW(5 *IW)) ff_ex_lpu_opc_bus (.CLK(clk), .LOAD(p_ce), .D(s1i_lpu_opc_bus), .Q(ex_lpu_opc_bus) );
   ysyx_20210479_mDFF_l # (.DW(8*IW)) ff_ex_epu_opc_bus (.CLK(clk), .LOAD(p_ce), .D(s1i_epu_opc_bus), .Q(ex_epu_opc_bus) );
   ysyx_20210479_mDFF_l # (.DW(8*IW)) ff_ex_bru_opc_bus (.CLK(clk), .LOAD(p_ce), .D(s1i_bru_opc_bus), .Q(ex_bru_opc_bus) );
   ysyx_20210479_mDFF_l # (.DW(7*IW)) ff_ex_lsu_opc_bus (.CLK(clk), .LOAD(p_ce), .D(s1i_lsu_opc_bus), .Q(ex_lsu_opc_bus) );
   ysyx_20210479_mDFF_l # (.DW((2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*IW)) ff_ex_bpu_upd (.CLK(clk), .LOAD(p_ce), .D(id_bpu_upd), .Q(ex_bpu_upd) );
   ysyx_20210479_mDFF_l # (.DW((CONFIG_AW-2 )*IW)) ff_ex_pc (.CLK(clk), .LOAD(p_ce), .D(id_pc), .Q(ex_pc) );
   ysyx_20210479_mDFF_l # (.DW(CONFIG_DW*IW)) ff_ex_imm (.CLK(clk), .LOAD(p_ce), .D(s1i_imm), .Q(ex_imm) );
   ysyx_20210479_mDFF_l # (.DW(IW)) ff_s1o_rf_rs2_re (.CLK(clk), .LOAD(p_ce), .D(rf_rs2_re), .Q(s1o_rf_rs2_re) );
   ysyx_20210479_mDFF_l # (.DW(IW)) ff_ex_rf_we (.CLK(clk), .LOAD(p_ce), .D(rf_we), .Q(ex_rf_we) );
   ysyx_20210479_mDFF_l # (.DW(5*IW)) ff_ex_rf_waddr (.CLK(clk), .LOAD(p_ce), .D(rf_waddr), .Q(ex_rf_waddr) );
endmodule
module ysyx_20210479_id_dec
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_ENABLE_MUL = 0,
   parameter                           CONFIG_ENABLE_DIV = 0,
   parameter                           CONFIG_ENABLE_DIVU = 0,
   parameter                           CONFIG_ENABLE_MOD = 0,
   parameter                           CONFIG_ENABLE_MODU = 0,
   parameter                           CONFIG_ENABLE_ASR = 0
)
(
   input                               id_valid,
   input [((2 <<1)*8)-1:0]           id_ins,
   input [2-1:0]              id_exc,
   input                               irq_async,
   output                              single_fu,
   output [9 -1:0]         alu_opc_bus,
   output [5 -1:0]         lpu_opc_bus,
   output [8-1:0]         epu_opc_bus,
   output [8-1:0]         bru_opc_bus,
   output [7-1:0]         lsu_opc_bus,
   output [CONFIG_DW-1:0]              imm,
   output                              rf_we,
   output [5-1:0]           rf_waddr,
   output                              rf_rs1_re,
   output [5-1:0]           rf_rs1_addr,
   output                              rf_rs2_re,
   output [5-1:0]           rf_rs2_addr
);
   wire                                msk;
   wire [6:0]                          f_opcode;
   wire [4:0]                          f_rd;
   wire [4:0]                          f_rs1;
   wire [4:0]                          f_rs2;
   wire [14:0]                         f_imm15;
   wire [16:0]                         f_imm17;
   wire [14:0]                         f_rel15;
   wire [24:0]                         f_rel25;
   wire                                enable_asr;
   wire                                enable_asr_i;
   wire                                enable_mul;
   wire                                enable_div;
   wire                                enable_divu;
   wire                                enable_mod;
   wire                                enable_modu;
   wire                                op_ldb;
   wire                                op_ldbu;
   wire                                op_ldh;
   wire                                op_ldhu;
   wire                                op_ldwu;
   wire                                op_stb;
   wire                                op_sth;
   wire                                op_stw;
   wire                                op_and;
   wire                                op_and_i;
   wire                                op_or;
   wire                                op_or_i;
   wire                                op_xor;
   wire                                op_xor_i;
   wire                                op_lsl;
   wire                                op_lsl_i;
   wire                                op_lsr;
   wire                                op_lsr_i;
   wire                                op_asr;
   wire                                op_asr_i;
   wire                                op_add;
   wire                                op_add_i;
   wire                                op_sub;
   wire                                op_mul;
   wire                                op_div;
   wire                                op_divu;
   wire                                op_mod;
   wire                                op_modu;
   wire                                op_mhi;
   wire                                op_jmp_i;
   wire                                op_jmp_lnk_i;
   wire                                op_jmpreg;
   wire                                op_beq;
   wire                                op_bne;
   wire                                op_bgt;
   wire                                op_bgtu;
   wire                                op_ble;
   wire                                op_bleu;
   wire                                op_syscall;
   wire                                op_ret;
   wire                                op_wmsr;
   wire                                op_rmsr;
   wire                                is_bcc;
   wire                                insn_rs1_imm15;
   wire                                insn_rd_rs1_imm15;
   wire                                insn_rd_rs1_rel15;
   wire                                insn_uimm17;
   wire                                insn_rel25;
   wire                                insn_no_rops;
   wire                                use_simm15;
   wire                                not_wb;
   wire                                read_rd_as_rs2;
   wire [CONFIG_DW-1:0]                imm15;
   wire [CONFIG_DW-1:0]                uimm17;
   wire [CONFIG_DW-1:0]                rel15;
   wire [CONFIG_DW-1:0]                rel25;
   wire [8-1:0]           epu_opc_no_EINSN;
   assign msk = ((~|id_exc) & ~irq_async & id_valid);
   assign f_opcode = id_ins[6:0] & {7{msk}}; 
   assign f_rd = id_ins[11:7];
   assign f_rs1 = id_ins[16:12];
   assign f_rs2 = id_ins[21:17];
   assign f_imm15 = id_ins[31:17];
   assign f_imm17 = id_ins[28:12];
   assign f_rel15 = id_ins[31:17];
   assign f_rel25 = id_ins[31:7];
   assign enable_asr = 1'b1;
   assign enable_asr_i = 1'b1;
   assign enable_mul = 1'b1;
   assign enable_div = 1'b1;
   assign enable_divu = 1'b1;
   assign enable_mod = 1'b1;
   assign enable_modu = 1'b1;
   assign op_ldb = (f_opcode == 7'h1d);
   assign op_ldbu = (f_opcode == 7'h1c);
   assign op_ldh = (f_opcode == 7'h1a);
   assign op_ldhu = (f_opcode == 7'h19);
   assign op_ldwu = (f_opcode == 7'h17);
   assign op_stb = (f_opcode == 7'h1e);
   assign op_sth = (f_opcode == 7'h1b);
   assign op_stw = (f_opcode == 7'h18);
   assign op_and = (f_opcode == 7'h0);
   assign op_and_i = (f_opcode == 7'h1);
   assign op_or = (f_opcode == 7'h2);
   assign op_or_i = (f_opcode == 7'h3);
   assign op_xor = (f_opcode == 7'h4);
   assign op_xor_i = (f_opcode == 7'h5);
   assign op_lsl = (f_opcode == 7'h6);
   assign op_lsl_i = (f_opcode == 7'h7);
   assign op_lsr = (f_opcode == 7'h8);
   assign op_lsr_i = (f_opcode == 7'h9);
   assign op_add = (f_opcode == 7'ha);
   assign op_add_i = (f_opcode == 7'hb);
   assign op_sub = (f_opcode == 7'hc);
   generate
      if (CONFIG_ENABLE_MUL)
         assign op_mul = (f_opcode == 7'h32) & enable_mul;
      else
         assign op_mul = 1'b0;
      if (CONFIG_ENABLE_DIV)
         assign op_div = (f_opcode == 7'h33) & enable_div;
      else
         assign op_div = 1'b0;
      if (CONFIG_ENABLE_DIVU)
         assign op_divu = (f_opcode == 7'h34) & enable_divu;
      else
         assign op_divu = 1'b0;
      if (CONFIG_ENABLE_MOD)
         assign op_mod = (f_opcode == 7'h35) & enable_mod;
      else
         assign op_mod = 1'b0;
      if (CONFIG_ENABLE_MODU)
         assign op_modu = (f_opcode == 7'h36) & enable_modu;
      else
         assign op_modu = 1'b0;
      if (CONFIG_ENABLE_ASR)
         begin
            assign op_asr = (f_opcode == 7'h30) & enable_asr;
            assign op_asr_i = (f_opcode == 7'h31) & enable_asr_i;
         end
      else
         begin
            assign op_asr = 1'b0;
            assign op_asr_i = 1'b0;
         end
   endgenerate
   assign op_mhi = (f_opcode == 7'h37);
   assign op_jmp_i = (f_opcode == 7'he);
   assign op_jmp_lnk_i = (f_opcode == 7'hf);
   assign op_jmpreg = (f_opcode == 7'hd);
   assign op_beq = (f_opcode == 7'h10);
   assign op_bne = (f_opcode == 7'h11);
   assign op_bgt = (f_opcode == 7'h12);
   assign op_bgtu = (f_opcode == 7'h13);
   assign op_ble = (f_opcode == 7'h14);
   assign op_bleu = (f_opcode == 7'h15);
   assign op_syscall = (f_opcode == 7'h21);
   assign op_ret = (f_opcode == 7'h22);
   assign op_wmsr = (f_opcode == 7'h23);
   assign op_rmsr = (f_opcode == 7'h24);
   assign alu_opc_bus[3] = (op_and | op_and_i);
   assign alu_opc_bus[4] = (op_or | op_or_i);
   assign alu_opc_bus[5] = (op_xor | op_xor_i);
   assign alu_opc_bus[6] = (op_lsl | op_lsl_i);
   assign alu_opc_bus[7] = (op_lsr | op_lsr_i);
   assign alu_opc_bus[8] = (op_asr | op_asr_i);
   assign alu_opc_bus[0] = (op_add | op_add_i);
   assign alu_opc_bus[1] = (op_sub);
   assign alu_opc_bus[2] = (op_mhi);
   assign bru_opc_bus[0] = (op_beq);
   assign bru_opc_bus[1] = (op_bne);
   assign bru_opc_bus[2] = (op_bgt);
   assign bru_opc_bus[3] = (op_bgtu);
   assign bru_opc_bus[4] = (op_ble);
   assign bru_opc_bus[5] = (op_bleu);
   assign bru_opc_bus[7] = (op_jmp_lnk_i | op_jmp_i);
   assign bru_opc_bus[6] = op_jmpreg;
   assign is_bcc = (op_beq | op_bne | op_bgt | op_bgtu | op_ble | op_bleu);
   assign lpu_opc_bus[0] = op_mul;
   assign lpu_opc_bus[1] = op_div;
   assign lpu_opc_bus[2] = op_divu;
   assign lpu_opc_bus[3] = op_mod;
   assign lpu_opc_bus[4] = op_modu;
   assign lsu_opc_bus[6:4] = (op_ldb|op_ldbu|op_stb)
                                          ? 3'd1
                                          : (op_ldh|op_ldhu|op_sth)
                                             ? 3'd2
                                             : (op_ldwu|op_stw)
                                                ? 3'd3
                                                : 3'd0;
   assign lsu_opc_bus[3] = (op_ldb | op_ldh);
   assign lsu_opc_bus[0] = (op_ldb|op_ldbu|op_ldh|op_ldhu|op_ldwu);
   assign lsu_opc_bus[1] = (op_stb|op_sth|op_stw);
   assign lsu_opc_bus[2] = (f_opcode == 7'h20);
   assign epu_opc_no_EINSN[0] = op_wmsr;
   assign epu_opc_no_EINSN[1] = op_rmsr;
   assign epu_opc_no_EINSN[2] = op_syscall;
   assign epu_opc_no_EINSN[3] = op_ret;
   assign epu_opc_no_EINSN[4] = (id_exc[0] & ~irq_async);
   assign epu_opc_no_EINSN[5] = (id_exc[1] & ~irq_async);
   assign epu_opc_no_EINSN[6] = irq_async;
   assign epu_opc_no_EINSN[(8-1)] = 1'b0;
   assign epu_opc_bus[(8-1)] =
      ~(
         (|alu_opc_bus) |
         (|lpu_opc_bus) |
         (|bru_opc_bus) |
         (lsu_opc_bus[0] | lsu_opc_bus[1] | lsu_opc_bus[2]) |
         (|epu_opc_no_EINSN)
      );
   assign epu_opc_bus[(8-1)-1:0] = epu_opc_no_EINSN[(8-1)-1:0];
   assign single_fu =
      (
         (|lpu_opc_bus) |
         (|bru_opc_bus) |
         (lsu_opc_bus[0] | lsu_opc_bus[1] | lsu_opc_bus[2]) |
         (|epu_opc_bus)
      );
   assign insn_rs1_imm15 =
      (
         op_and_i | op_or_i | op_xor_i | op_lsl_i | op_lsr_i | op_asr_i |
         op_add_i |
         lsu_opc_bus[0] |
         op_rmsr
      );
   assign insn_rd_rs1_imm15 =
      (
         lsu_opc_bus[1] |
         op_wmsr
      );
   assign insn_rd_rs1_rel15 = is_bcc;
   assign insn_uimm17 = op_mhi;
   assign insn_rel25 = (op_jmp_i | op_jmp_lnk_i);
   assign use_simm15 = (op_xor_i | op_add_i | lsu_opc_bus[0] | lsu_opc_bus[1]);
   assign insn_no_rops = (op_mhi | lsu_opc_bus[2] | op_syscall | op_ret | op_jmp_i | op_jmp_lnk_i);
   assign not_wb =
      (
         op_jmp_i | is_bcc | 
         lsu_opc_bus[1] | lsu_opc_bus[2] |
         op_wmsr | epu_opc_bus[2] | epu_opc_bus[3] |
         epu_opc_bus[4] | epu_opc_bus[5] |
         epu_opc_bus[(8-1)] |
         epu_opc_bus[6]
      );
   assign rf_we = ~not_wb & (|rf_waddr);
   assign rf_waddr = (op_jmp_lnk_i) ? 1  : f_rd;
   assign read_rd_as_rs2 = (lsu_opc_bus[1] | op_wmsr | is_bcc);
   assign rf_rs1_re = ~insn_no_rops;
   assign rf_rs1_addr = f_rs1;
   assign rf_rs2_re = ((~insn_rs1_imm15 & ~insn_uimm17 & ~insn_rel25 & ~insn_no_rops) | read_rd_as_rs2);
   assign rf_rs2_addr = read_rd_as_rs2 ? f_rd : f_rs2;
   assign imm15 = {{CONFIG_DW-15{use_simm15 & f_imm15[14]}}, f_imm15[14:0]};
   assign uimm17 = {{CONFIG_DW-17{1'b0}}, f_imm17[16:0]};
   assign rel15 = {{CONFIG_DW-2-15{f_rel15[14]}}, f_rel15[14:0], 2'b00};
   assign rel25 = {{CONFIG_DW-2-25{f_rel25[24]}}, f_rel25[24:0], 2'b00};
   assign imm = ({CONFIG_DW{insn_rs1_imm15|insn_rd_rs1_imm15}} & imm15) |
                  ({CONFIG_DW{insn_rd_rs1_rel15}} & rel15) |
                  ({CONFIG_DW{insn_rel25}} & rel25) |
                  ({CONFIG_DW{insn_uimm17}} & uimm17);
endmodule
module ysyx_20210479_id_ro
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_P_ISSUE_WIDTH = 0
)
(
   input                               clk,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_dout,
   input [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_wdat,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_we,
   input [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_we,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_waddr,
   input [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_waddr,
   input ro_ex_s1_load0,
   input ro_ex_s2_load0,
   input ro_ex_s3_load0,
   input [5*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] raddr,
   input [2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] re,
   input [CONFIG_DW*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] rf_din,
   output [CONFIG_DW*2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] byp_dout,
   output [2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] raw_dep_load0
);
   localparam IW                       = (1<<CONFIG_P_ISSUE_WIDTH);
   localparam CHS                      = (IW*2);
   wire                                p_ce;
   wire [CONFIG_DW*IW-1:0]             s1o_ex_s1_rf_dout_ff, s1o_ex_s1_rf_dout_ff_rev;
   wire [CONFIG_DW*IW-1:0]             s1o_ex_s2_rf_dout_ff, s1o_ex_s2_rf_dout_ff_rev;
   wire [CONFIG_DW*IW-1:0]             s1o_ex_s3_rf_dout_ff, s1o_ex_s3_rf_dout_ff_rev;
   wire [CONFIG_DW*IW-1:0]             s1o_cmt_rf_wdat_ff, s1o_cmt_rf_wdat_ff_rev;
   wire [CHS-1:0]                      rop_raw_load0;
   genvar i, k;
   integer j;
   generate
      for(i=0;i<CHS;i=i+1)
         begin
            wire [IW-1:0]        cf_ex_s1, cf_ex_s2, cf_ex_s3, cf_cmt;
            wire [IW-1:0]        cf_ex_s1_rev, cf_ex_s2_rev, cf_ex_s3_rev, cf_cmt_rev;
            wire [IW-1:0]        s1o_cf_ex_s1_rev, s1o_cf_ex_s2_rev, s1o_cf_ex_s3_rev, s1o_cf_cmt_rev;
            wire                 s1o_use_ex_s1, s1o_use_ex_s2, s1o_use_ex_s3, s1o_use_cmt;
            wire [CONFIG_DW-1:0] s1o_ex_s1_rf_dout_sel;
            wire [CONFIG_DW-1:0] s1o_ex_s2_rf_dout_sel;
            wire [CONFIG_DW-1:0] s1o_ex_s3_rf_dout_sel;
            wire [CONFIG_DW-1:0] s1o_cmt_rf_wdat_sel;
            for(k=0;k<IW;k=k+1)
               begin
                  assign cf_ex_s1[k] = ((raddr[i*5 +: 5] == ro_ex_s1_rf_waddr[k*5 +: 5]) &
                                       re[i] & ro_ex_s1_rf_we[k]);
                  assign cf_ex_s2[k] = ((raddr[i*5 +: 5] == ro_ex_s2_rf_waddr[k*5 +: 5]) &
                                       re[i] & ro_ex_s2_rf_we[k]);
                  assign cf_ex_s3[k] = ((raddr[i*5 +: 5] == ro_ex_s3_rf_waddr[k*5 +: 5]) &
                                       re[i] & ro_ex_s3_rf_we[k]);
                  assign cf_cmt[k] = ((raddr[i*5 +: 5] == ro_cmt_rf_waddr[k*5 +: 5]) &
                                       re[i] & ro_cmt_rf_we[k]);
                  assign cf_ex_s1_rev[IW-k-1] = cf_ex_s1[k];
                  assign cf_ex_s2_rev[IW-k-1] = cf_ex_s2[k];
                  assign cf_ex_s3_rev[IW-k-1] = cf_ex_s3[k];
                  assign cf_cmt_rev[IW-k-1] = cf_cmt[k];
               end
            assign raw_dep_load0[i] = (cf_ex_s1[0] & ro_ex_s1_load0) |
                                       (cf_ex_s2[0] & ro_ex_s2_load0) |
                                       (cf_ex_s3[0] & ro_ex_s3_load0);
            ysyx_20210479_mDFF_l #(.DW(IW)) ff_s1o_cf_ex_s1_rev(.CLK(clk), .LOAD(p_ce), .D(cf_ex_s1_rev), .Q(s1o_cf_ex_s1_rev) );
            ysyx_20210479_mDFF_l #(.DW(IW)) ff_s1o_cf_ex_s2_rev(.CLK(clk), .LOAD(p_ce), .D(cf_ex_s2_rev), .Q(s1o_cf_ex_s2_rev) );
            ysyx_20210479_mDFF_l #(.DW(IW)) ff_s1o_cf_ex_s3_rev(.CLK(clk), .LOAD(p_ce), .D(cf_ex_s3_rev), .Q(s1o_cf_ex_s3_rev) );
            ysyx_20210479_mDFF_l #(.DW(IW)) ff_s1o_cf_cmt_rev(.CLK(clk), .LOAD(p_ce), .D(cf_cmt_rev), .Q(s1o_cf_cmt_rev) );
            ysyx_20210479_pmux_v #(.SELW(IW), .DW(CONFIG_DW)) U_EX_S1_PMUX (.sel(s1o_cf_ex_s1_rev), .din(s1o_ex_s1_rf_dout_ff_rev), .dout(s1o_ex_s1_rf_dout_sel), .valid(s1o_use_ex_s1) );
            ysyx_20210479_pmux_v #(.SELW(IW), .DW(CONFIG_DW)) U_EX_S2_PMUX (.sel(s1o_cf_ex_s2_rev), .din(s1o_ex_s2_rf_dout_ff_rev), .dout(s1o_ex_s2_rf_dout_sel), .valid(s1o_use_ex_s2) );
            ysyx_20210479_pmux_v #(.SELW(IW), .DW(CONFIG_DW)) U_EX_S3_PMUX (.sel(s1o_cf_ex_s3_rev), .din(s1o_ex_s3_rf_dout_ff_rev), .dout(s1o_ex_s3_rf_dout_sel), .valid(s1o_use_ex_s3) );
            ysyx_20210479_pmux_v #(.SELW(IW), .DW(CONFIG_DW)) U_CMT_PMUX (.sel(s1o_cf_cmt_rev), .din(s1o_cmt_rf_wdat_ff_rev), .dout(s1o_cmt_rf_wdat_sel), .valid(s1o_use_cmt) );
            assign byp_dout[i*CONFIG_DW +: CONFIG_DW] = (s1o_use_ex_s1)
                                                            ? s1o_ex_s1_rf_dout_sel
                                                            : (s1o_use_ex_s2)
                                                               ? s1o_ex_s2_rf_dout_sel
                                                               : (s1o_use_ex_s3)
                                                                  ? s1o_ex_s3_rf_dout_sel
                                                                  : (s1o_use_cmt)
                                                                     ? s1o_cmt_rf_wdat_sel
                                                                     : rf_din[i*CONFIG_DW +: CONFIG_DW];
         end
   endgenerate
   assign p_ce = (|re);
   ysyx_20210479_mDFF_l #(.DW(CONFIG_DW*IW)) ff_s1o_ex_s1_rf_dout_ff(.CLK(clk), .LOAD(p_ce), .D(ro_ex_s1_rf_dout), .Q(s1o_ex_s1_rf_dout_ff) );
   ysyx_20210479_mDFF_l #(.DW(CONFIG_DW*IW)) ff_s1o_ex_s2_rf_dout_ff(.CLK(clk), .LOAD(p_ce), .D(ro_ex_s2_rf_dout), .Q(s1o_ex_s2_rf_dout_ff) );
   ysyx_20210479_mDFF_l #(.DW(CONFIG_DW*IW)) ff_s1o_ex_s3_rf_wdat_ff(.CLK(clk), .LOAD(p_ce), .D(ro_ex_s3_rf_dout), .Q(s1o_ex_s3_rf_dout_ff) );
   ysyx_20210479_mDFF_l #(.DW(CONFIG_DW*IW)) ff_s1o_cmt_rf_wdat_ff(.CLK(clk), .LOAD(p_ce), .D(ro_cmt_rf_wdat), .Q(s1o_cmt_rf_wdat_ff) );
   generate
      for(i=0;i<IW;i=i+1)
         begin : gen_s1o_rf_dout_ff_rev
            assign s1o_ex_s1_rf_dout_ff_rev[(IW-i-1)*CONFIG_DW +: CONFIG_DW] = s1o_ex_s1_rf_dout_ff[i*CONFIG_DW +: CONFIG_DW];
            assign s1o_ex_s2_rf_dout_ff_rev[(IW-i-1)*CONFIG_DW +: CONFIG_DW] = s1o_ex_s2_rf_dout_ff[i*CONFIG_DW +: CONFIG_DW];
            assign s1o_ex_s3_rf_dout_ff_rev[(IW-i-1)*CONFIG_DW +: CONFIG_DW] = s1o_ex_s3_rf_dout_ff[i*CONFIG_DW +: CONFIG_DW];
            assign s1o_cmt_rf_wdat_ff_rev[(IW-i-1)*CONFIG_DW +: CONFIG_DW] = s1o_cmt_rf_wdat_ff[i*CONFIG_DW +: CONFIG_DW];
         end
   endgenerate
endmodule
module ysyx_20210479_immu
#(
   parameter                           CONFIG_AW = 0,
   parameter                           CONFIG_DW = 0,
   parameter                           CONFIG_IMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_P_PAGE_SIZE = 0,
   parameter                           CONFIG_ITLB_P_SETS = 0
)
(
   input                               clk,
   input                               rst,
   input                               re,
   input [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] vpn,
   output [CONFIG_AW-CONFIG_P_PAGE_SIZE-1:0] ppn,
   output                              EITM,
   output                              EIPF,
   output                              uncached,
   input                               msr_psr_imme,
   input                               msr_psr_rm,
   output [CONFIG_DW-1:0]              msr_immid,
   input [CONFIG_ITLB_P_SETS-1:0]      msr_imm_tlbl_idx,
   input [CONFIG_DW-1:0]               msr_imm_tlbl_nxt,
   input                               msr_imm_tlbl_we,
   input [CONFIG_ITLB_P_SETS-1:0]      msr_imm_tlbh_idx,
   input [CONFIG_DW-1:0]               msr_imm_tlbh_nxt,
   input                               msr_imm_tlbh_we
);
   localparam VPN_SHIFT                = CONFIG_P_PAGE_SIZE;
   localparam PPN_SHIFT                = VPN_SHIFT;
   localparam VPN_DW                   = CONFIG_AW-VPN_SHIFT;
   localparam PPN_DW                   = CONFIG_AW-PPN_SHIFT;
   assign msr_immid = {{32-3{1'b0}}, CONFIG_ITLB_P_SETS[2:0]};
   wire                                msr_psr_imme_ff;
   wire                                msr_psr_rm_ff;
   wire [VPN_DW-1:0]                   tgt_vpn_ff;
   wire [CONFIG_DW-1:0]                tlb_l_ff;
   wire [CONFIG_DW-1:0]                tlb_h_ff;
   wire [VPN_DW-1:0] tgt_vpn_nxt = vpn[VPN_DW-1:0];
   wire [CONFIG_ITLB_P_SETS-1:0] tgt_index_nxt = tgt_vpn_nxt[CONFIG_ITLB_P_SETS-1:0];
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_imme (.CLK(clk),.RST(rst), .LOAD(re), .D(msr_psr_imme), .Q(msr_psr_imme_ff) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_msr_psr_rm (.CLK(clk),.RST(rst), .LOAD(re), .D(msr_psr_rm), .Q(msr_psr_rm_ff) );
   ysyx_20210479_mDFF_lr #(.DW(VPN_DW)) ff_tgt_vpn (.CLK(clk),.RST(rst), .LOAD(re), .D(tgt_vpn_nxt), .Q(tgt_vpn_ff) );
   ysyx_20210479_mRF_nwnr
      #(
         .DW      (CONFIG_DW),
         .AW      (CONFIG_ITLB_P_SETS),
         .NUM_READ (1),
         .NUM_WRITE (1)
      )
   U_TLB_L
      (
         .CLK     (clk),
         .RE      (re),
         .RADDR   (tgt_index_nxt),
         .RDATA   (tlb_l_ff),
         .WE      (msr_imm_tlbl_we),
         .WADDR   (msr_imm_tlbl_idx),
         .WDATA   (msr_imm_tlbl_nxt)
      );
   ysyx_20210479_mRF_nwnr
      #(
         .DW      (CONFIG_DW),
         .AW      (CONFIG_ITLB_P_SETS),
         .NUM_READ (1),
         .NUM_WRITE (1)
      )
   U_TLB_H
      (
         .CLK     (clk),
         .RE      (re),
         .RADDR   (tgt_index_nxt),
         .RDATA   (tlb_h_ff),
         .WE      (msr_imm_tlbh_we),
         .WADDR   (msr_imm_tlbh_idx),
         .WDATA   (msr_imm_tlbh_nxt)
      );
   wire tlb_v = tlb_l_ff[0];
   wire [VPN_DW-1:0] tlb_vpn = tlb_l_ff[CONFIG_DW-1:CONFIG_DW-VPN_DW];
   wire tlb_p = tlb_h_ff[0];
   wire tlb_ux = tlb_h_ff[3];
   wire tlb_rx = tlb_h_ff[4];
   wire tlb_unc = tlb_h_ff[7];
   wire tlb_s = tlb_h_ff[8];
   wire [PPN_DW-1:0] tlb_ppn = tlb_h_ff[CONFIG_DW-1:CONFIG_DW-PPN_DW];
   wire perm_denied;
   wire tlb_miss;
   assign perm_denied =
      (
         (msr_psr_rm_ff & ~tlb_rx) |
         (~msr_psr_rm_ff & ~tlb_ux)
      );
   assign tlb_miss = ~(tlb_v & tlb_vpn == tgt_vpn_ff);
   assign EITM = (tlb_miss & msr_psr_imme_ff);
   assign EIPF = (perm_denied & ~tlb_miss & msr_psr_imme_ff);
   assign ppn = msr_psr_imme_ff ? tlb_ppn : tgt_vpn_ff;
generate
   if (CONFIG_IMMU_ENABLE_UNCACHED_SEG)
      assign uncached = (msr_psr_imme_ff & ~tlb_miss & ~perm_denied & tlb_unc) | (~EITM & ~EIPF & ~ppn[CONFIG_AW-CONFIG_P_PAGE_SIZE-1]);
   else
      assign uncached = (msr_psr_imme_ff & ~tlb_miss & ~perm_denied & tlb_unc);
endgenerate
endmodule
module ysyx_20210479_ncpu64k
#(
   parameter                           CONFIG_AW = 32,
   parameter                           CONFIG_DW = 32,
   parameter                           CONFIG_P_DW = 5,
   parameter                           CONFIG_P_FETCH_WIDTH = 1,
   parameter                           CONFIG_P_ISSUE_WIDTH = 1,
   parameter                           CONFIG_P_PAGE_SIZE = 13,
   parameter                           CONFIG_IC_P_LINE = 6,
   parameter                           CONFIG_IC_P_SETS = 6,
   parameter                           CONFIG_IC_P_WAYS = 2,
   parameter                           CONFIG_DC_P_LINE = 6,
   parameter                           CONFIG_DC_P_SETS = 6,
   parameter                           CONFIG_DC_P_WAYS = 2,
   parameter                           CONFIG_PHT_P_NUM = 9,
   parameter                           CONFIG_BTB_P_NUM = 9,
   parameter                           CONFIG_P_IQ_DEPTH = 4,
   parameter                           CONFIG_ENABLE_MUL = 0,
   parameter                           CONFIG_ENABLE_DIV = 0,
   parameter                           CONFIG_ENABLE_DIVU = 0,
   parameter                           CONFIG_ENABLE_MOD = 0,
   parameter                           CONFIG_ENABLE_MODU = 0,
   parameter                           CONFIG_ENABLE_ASR = 0,
   parameter                           CONFIG_IMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_DMMU_ENABLE_UNCACHED_SEG = 0,
   parameter                           CONFIG_DTLB_P_SETS = 7,
   parameter                           CONFIG_ITLB_P_SETS = 7,
   parameter [CONFIG_AW-1:0]           CONFIG_ERST_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EITM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_ESYSCALL_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EINSN_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EIRQ_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDTM_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EDPF_VECTOR = 0,
   parameter [CONFIG_AW-1:0]           CONFIG_EALIGN_VECTOR = 0,
   parameter                           CONFIG_NUM_IRQ = 32,
   parameter                           AXI_P_DW_BYTES    = 3,
   parameter                           AXI_UNCACHED_P_DW_BYTES = 2,
   parameter                           AXI_ADDR_WIDTH    = 64,
   parameter                           AXI_ID_WIDTH      = 4,
   parameter                           AXI_USER_WIDTH    = 1
)
(
   input                               clk,
   input                               rst,
   input                               ibus_ARREADY,
   output                              ibus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         ibus_ARADDR,
   output [2:0]                        ibus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           ibus_ARID,
   output [AXI_USER_WIDTH-1:0]         ibus_ARUSER,
   output [7:0]                        ibus_ARLEN,
   output [2:0]                        ibus_ARSIZE,
   output [1:0]                        ibus_ARBURST,
   output                              ibus_ARLOCK,
   output [3:0]                        ibus_ARCACHE,
   output [3:0]                        ibus_ARQOS,
   output [3:0]                        ibus_ARREGION,
   output                              ibus_RREADY,
   input                               ibus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  ibus_RDATA,
   input                               ibus_RLAST,
   input  [1:0]                        ibus_RRESP,
   input  [AXI_ID_WIDTH-1:0]           ibus_RID,
   input  [AXI_USER_WIDTH-1:0]         ibus_RUSER,
   input                               dbus_ARREADY,
   output                              dbus_ARVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_ARADDR,
   output [2:0]                        dbus_ARPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_ARID,
   output [AXI_USER_WIDTH-1:0]         dbus_ARUSER,
   output [7:0]                        dbus_ARLEN,
   output [2:0]                        dbus_ARSIZE,
   output [1:0]                        dbus_ARBURST,
   output                              dbus_ARLOCK,
   output [3:0]                        dbus_ARCACHE,
   output [3:0]                        dbus_ARQOS,
   output [3:0]                        dbus_ARREGION,
   output                              dbus_RREADY,
   input                               dbus_RVALID,
   input  [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_RDATA,
   input  [1:0]                        dbus_RRESP,
   input                               dbus_RLAST,
   input  [AXI_ID_WIDTH-1:0]           dbus_RID,
   input  [AXI_USER_WIDTH-1:0]         dbus_RUSER,
   input                               dbus_AWREADY,
   output                              dbus_AWVALID,
   output [AXI_ADDR_WIDTH-1:0]         dbus_AWADDR,
   output [2:0]                        dbus_AWPROT,
   output [AXI_ID_WIDTH-1:0]           dbus_AWID,
   output [AXI_USER_WIDTH-1:0]         dbus_AWUSER,
   output [7:0]                        dbus_AWLEN,
   output [2:0]                        dbus_AWSIZE,
   output [1:0]                        dbus_AWBURST,
   output                              dbus_AWLOCK,
   output [3:0]                        dbus_AWCACHE,
   output [3:0]                        dbus_AWQOS,
   output [3:0]                        dbus_AWREGION,
   input                               dbus_WREADY,
   output                              dbus_WVALID,
   output [(1<<AXI_P_DW_BYTES)*8-1:0]  dbus_WDATA,
   output [(1<<AXI_P_DW_BYTES)-1:0]    dbus_WSTRB,
   output                              dbus_WLAST,
   output [AXI_USER_WIDTH-1:0]         dbus_WUSER,
   output                              dbus_BREADY,
   input                               dbus_BVALID,
   input [1:0]                         dbus_BRESP,
   input [AXI_ID_WIDTH-1:0]            dbus_BID,
   input [AXI_USER_WIDTH-1:0]          dbus_BUSER,
   input [CONFIG_NUM_IRQ-1:0]          irqs,
   output                              tsc_irq
);
   wire [(1<<CONFIG_P_ISSUE_WIDTH)*2*5-1:0] arf_RADDR;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)*2*CONFIG_DW-1:0] arf_RDATA;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)*2-1:0] arf_RE;
   wire                 bpu_wb;                 
   wire                 bpu_wb_is_bcc;          
   wire                 bpu_wb_is_breg;         
   wire                 bpu_wb_is_brel;         
   wire [(CONFIG_AW-2 )-1:0]     bpu_wb_npc_act;         
   wire [(CONFIG_AW-2 )-1:0]     bpu_wb_pc;              
   wire                 bpu_wb_taken;           
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0] bpu_wb_upd;            
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_waddr;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_wdat;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] commit_rf_we;
   wire [9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_alu_opc_bus;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bpu_upd;
   wire [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_bru_opc_bus;
   wire [8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_epu_opc_bus;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_imm;
   wire [5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lpu_opc_bus;
   wire [7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_lsu_opc_bus;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand1;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_operand2;
   wire [(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_pc;
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_waddr;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_rf_we;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ex_valid;
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_bpu_upd;
   wire [2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_exc;
   wire [((2 <<1)*8)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_ins;
   wire [(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_pc;
   wire [CONFIG_P_ISSUE_WIDTH:0] id_pop_cnt;    
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_valid;
   wire                 irq_async;              
   wire [CONFIG_DW-1:0] msr_icid;               
   wire [CONFIG_DW-1:0] msr_icinv_nxt;          
   wire                 msr_icinv_ready;        
   wire                 msr_icinv_we;           
   wire [CONFIG_ITLB_P_SETS-1:0] msr_imm_tlbh_idx;
   wire [CONFIG_DW-1:0] msr_imm_tlbh_nxt;       
   wire                 msr_imm_tlbh_we;        
   wire [CONFIG_ITLB_P_SETS-1:0] msr_imm_tlbl_idx;
   wire [CONFIG_DW-1:0] msr_imm_tlbl_nxt;       
   wire                 msr_imm_tlbl_we;        
   wire [CONFIG_DW-1:0] msr_immid;              
   wire                 msr_psr_ice;            
   wire                 msr_psr_imme;           
   wire                 msr_psr_rm;             
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_waddr;
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_wdat;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_cmt_rf_we;
   wire                 ro_ex_s1_load0;         
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_dout;
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_waddr;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s1_rf_we;
   wire                 ro_ex_s2_load0;         
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_dout;
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_waddr;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s2_rf_we;
   wire                 ro_ex_s3_load0;         
   wire [CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_dout;
   wire [5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_waddr;
   wire [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] ro_ex_s3_rf_we;
   wire                                flush;                  
   wire [(CONFIG_AW-2 )-1:0]                    flush_tgt;             
   wire                                stall;                  
   ysyx_20210479_frontend
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH),
        .CONFIG_P_IQ_DEPTH              (CONFIG_P_IQ_DEPTH),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_ITLB_P_SETS             (CONFIG_ITLB_P_SETS),
        .CONFIG_IC_P_LINE               (CONFIG_IC_P_LINE),
        .CONFIG_IC_P_SETS               (CONFIG_IC_P_SETS),
        .CONFIG_IC_P_WAYS               (CONFIG_IC_P_WAYS),
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_ERST_VECTOR             (CONFIG_ERST_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_IMMU_ENABLE_UNCACHED_SEG(CONFIG_IMMU_ENABLE_UNCACHED_SEG),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_UNCACHED_P_DW_BYTES        (AXI_UNCACHED_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_FNT
      (
       .id_valid                        (id_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_ins                          (id_ins[((2 <<1)*8)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_pc                           (id_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_exc                          (id_exc[2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_bpu_upd                      (id_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .msr_immid                       (msr_immid[CONFIG_DW-1:0]),
       .msr_icid                        (msr_icid[CONFIG_DW-1:0]),
       .msr_icinv_ready                 (msr_icinv_ready),
       .ibus_ARVALID                    (ibus_ARVALID),
       .ibus_ARADDR                     (ibus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .ibus_ARPROT                     (ibus_ARPROT[2:0]),
       .ibus_ARID                       (ibus_ARID[AXI_ID_WIDTH-1:0]),
       .ibus_ARUSER                     (ibus_ARUSER[AXI_USER_WIDTH-1:0]),
       .ibus_ARLEN                      (ibus_ARLEN[7:0]),
       .ibus_ARSIZE                     (ibus_ARSIZE[2:0]),
       .ibus_ARBURST                    (ibus_ARBURST[1:0]),
       .ibus_ARLOCK                     (ibus_ARLOCK),
       .ibus_ARCACHE                    (ibus_ARCACHE[3:0]),
       .ibus_ARQOS                      (ibus_ARQOS[3:0]),
       .ibus_ARREGION                   (ibus_ARREGION[3:0]),
       .ibus_RREADY                     (ibus_RREADY),
       .clk                             (clk),
       .rst                             (rst),
       .flush                           (flush),
       .flush_tgt                       (flush_tgt[(CONFIG_AW-2 )-1:0]),
       .id_pop_cnt                      (id_pop_cnt[CONFIG_P_ISSUE_WIDTH:0]),
       .bpu_wb                          (bpu_wb),
       .bpu_wb_is_bcc                   (bpu_wb_is_bcc),
       .bpu_wb_is_breg                  (bpu_wb_is_breg),
       .bpu_wb_is_brel                  (bpu_wb_is_brel),
       .bpu_wb_taken                    (bpu_wb_taken),
       .bpu_wb_pc                       (bpu_wb_pc[(CONFIG_AW-2 )-1:0]),
       .bpu_wb_npc_act                  (bpu_wb_npc_act[(CONFIG_AW-2 )-1:0]),
       .bpu_wb_upd                      (bpu_wb_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]),
       .msr_psr_imme                    (msr_psr_imme),
       .msr_psr_rm                      (msr_psr_rm),
       .msr_psr_ice                     (msr_psr_ice),
       .msr_imm_tlbl_idx                (msr_imm_tlbl_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbl_nxt                (msr_imm_tlbl_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbl_we                 (msr_imm_tlbl_we),
       .msr_imm_tlbh_idx                (msr_imm_tlbh_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbh_nxt                (msr_imm_tlbh_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbh_we                 (msr_imm_tlbh_we),
       .msr_icinv_nxt                   (msr_icinv_nxt[CONFIG_DW-1:0]),
       .msr_icinv_we                    (msr_icinv_we),
       .ibus_ARREADY                    (ibus_ARREADY),
       .ibus_RVALID                     (ibus_RVALID),
       .ibus_RDATA                      (ibus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .ibus_RRESP                      (ibus_RRESP[1:0]),
       .ibus_RLAST                      (ibus_RLAST),
       .ibus_RID                        (ibus_RID[AXI_ID_WIDTH-1:0]),
       .ibus_RUSER                      (ibus_RUSER[AXI_USER_WIDTH-1:0]));
   ysyx_20210479_id
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH),
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_ENABLE_MUL              (CONFIG_ENABLE_MUL),
        .CONFIG_ENABLE_DIV              (CONFIG_ENABLE_DIV),
        .CONFIG_ENABLE_DIVU             (CONFIG_ENABLE_DIVU),
        .CONFIG_ENABLE_MOD              (CONFIG_ENABLE_MOD),
        .CONFIG_ENABLE_MODU             (CONFIG_ENABLE_MODU),
        .CONFIG_ENABLE_ASR              (CONFIG_ENABLE_ASR))
   U_ID
      (
       .id_pop_cnt                      (id_pop_cnt[CONFIG_P_ISSUE_WIDTH:0]),
       .ex_valid                        (ex_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_alu_opc_bus                  (ex_alu_opc_bus[9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_lpu_opc_bus                  (ex_lpu_opc_bus[5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_epu_opc_bus                  (ex_epu_opc_bus[8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_bru_opc_bus                  (ex_bru_opc_bus[8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_lsu_opc_bus                  (ex_lsu_opc_bus[7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_bpu_upd                      (ex_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_pc                           (ex_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_imm                          (ex_imm[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_operand1                     (ex_operand1[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_operand2                     (ex_operand2[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_rf_waddr                     (ex_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_rf_we                        (ex_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .arf_RE                          (arf_RE[(1<<CONFIG_P_ISSUE_WIDTH)*2-1:0]),
       .arf_RADDR                       (arf_RADDR[(1<<CONFIG_P_ISSUE_WIDTH)*2*5-1:0]),
       .clk                             (clk),
       .rst                             (rst),
       .flush                           (flush),
       .stall                           (stall),
       .id_valid                        (id_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_ins                          (id_ins[((2 <<1)*8)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_pc                           (id_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_exc                          (id_exc[2*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .id_bpu_upd                      (id_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .irq_async                       (irq_async),
       .ro_ex_s1_rf_dout                (ro_ex_s1_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_dout                (ro_ex_s2_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_dout                (ro_ex_s3_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_wdat                  (ro_cmt_rf_wdat[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_we                  (ro_ex_s1_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_we                  (ro_ex_s2_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_we                  (ro_ex_s3_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_we                    (ro_cmt_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_waddr               (ro_ex_s1_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_waddr               (ro_ex_s2_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_waddr               (ro_ex_s3_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_waddr                 (ro_cmt_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_load0                  (ro_ex_s1_load0),
       .ro_ex_s2_load0                  (ro_ex_s2_load0),
       .ro_ex_s3_load0                  (ro_ex_s3_load0),
       .arf_RDATA                       (arf_RDATA[(1<<CONFIG_P_ISSUE_WIDTH)*2*CONFIG_DW-1:0]));
   ysyx_20210479_ex
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_DW                    (CONFIG_P_DW),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH),
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_ENABLE_MUL              (CONFIG_ENABLE_MUL),
        .CONFIG_ENABLE_DIV              (CONFIG_ENABLE_DIV),
        .CONFIG_ENABLE_DIVU             (CONFIG_ENABLE_DIVU),
        .CONFIG_ENABLE_MOD              (CONFIG_ENABLE_MOD),
        .CONFIG_ENABLE_MODU             (CONFIG_ENABLE_MODU),
        .CONFIG_ENABLE_ASR              (CONFIG_ENABLE_ASR),
        .CONFIG_NUM_IRQ                 (CONFIG_NUM_IRQ),
        .CONFIG_DC_P_WAYS               (CONFIG_DC_P_WAYS),
        .CONFIG_DC_P_SETS               (CONFIG_DC_P_SETS),
        .CONFIG_DC_P_LINE               (CONFIG_DC_P_LINE),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_DMMU_ENABLE_UNCACHED_SEG(CONFIG_DMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_ITLB_P_SETS             (CONFIG_ITLB_P_SETS),
        .CONFIG_DTLB_P_SETS             (CONFIG_DTLB_P_SETS),
        .CONFIG_EITM_VECTOR             (CONFIG_EITM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIPF_VECTOR             (CONFIG_EIPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_ESYSCALL_VECTOR         (CONFIG_ESYSCALL_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EINSN_VECTOR            (CONFIG_EINSN_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIRQ_VECTOR             (CONFIG_EIRQ_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDTM_VECTOR             (CONFIG_EDTM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDPF_VECTOR             (CONFIG_EDPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EALIGN_VECTOR           (CONFIG_EALIGN_VECTOR[CONFIG_AW-1:0]),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_EX
      (
       .stall                           (stall),
       .flush                           (flush),
       .flush_tgt                       (flush_tgt[(CONFIG_AW-2 )-1:0]),
       .ro_ex_s1_rf_dout                (ro_ex_s1_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_dout                (ro_ex_s2_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_dout                (ro_ex_s3_rf_dout[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_wdat                  (ro_cmt_rf_wdat[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_we                  (ro_ex_s1_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_we                  (ro_ex_s2_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_we                  (ro_ex_s3_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_we                    (ro_cmt_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_rf_waddr               (ro_ex_s1_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s2_rf_waddr               (ro_ex_s2_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s3_rf_waddr               (ro_ex_s3_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_cmt_rf_waddr                 (ro_cmt_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ro_ex_s1_load0                  (ro_ex_s1_load0),
       .ro_ex_s2_load0                  (ro_ex_s2_load0),
       .ro_ex_s3_load0                  (ro_ex_s3_load0),
       .commit_rf_wdat                  (commit_rf_wdat[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .commit_rf_waddr                 (commit_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .commit_rf_we                    (commit_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .bpu_wb                          (bpu_wb),
       .bpu_wb_is_bcc                   (bpu_wb_is_bcc),
       .bpu_wb_is_breg                  (bpu_wb_is_breg),
       .bpu_wb_is_brel                  (bpu_wb_is_brel),
       .bpu_wb_taken                    (bpu_wb_taken),
       .bpu_wb_pc                       (bpu_wb_pc[(CONFIG_AW-2 )-1:0]),
       .bpu_wb_npc_act                  (bpu_wb_npc_act[(CONFIG_AW-2 )-1:0]),
       .bpu_wb_upd                      (bpu_wb_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]),
       .irq_async                       (irq_async),
       .tsc_irq                         (tsc_irq),
       .msr_psr_imme                    (msr_psr_imme),
       .msr_psr_rm                      (msr_psr_rm),
       .msr_psr_ice                     (msr_psr_ice),
       .msr_imm_tlbl_idx                (msr_imm_tlbl_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbl_nxt                (msr_imm_tlbl_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbl_we                 (msr_imm_tlbl_we),
       .msr_imm_tlbh_idx                (msr_imm_tlbh_idx[CONFIG_ITLB_P_SETS-1:0]),
       .msr_imm_tlbh_nxt                (msr_imm_tlbh_nxt[CONFIG_DW-1:0]),
       .msr_imm_tlbh_we                 (msr_imm_tlbh_we),
       .msr_icinv_nxt                   (msr_icinv_nxt[CONFIG_DW-1:0]),
       .msr_icinv_we                    (msr_icinv_we),
       .dbus_ARVALID                    (dbus_ARVALID),
       .dbus_ARADDR                     (dbus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_ARPROT                     (dbus_ARPROT[2:0]),
       .dbus_ARID                       (dbus_ARID[AXI_ID_WIDTH-1:0]),
       .dbus_ARUSER                     (dbus_ARUSER[AXI_USER_WIDTH-1:0]),
       .dbus_ARLEN                      (dbus_ARLEN[7:0]),
       .dbus_ARSIZE                     (dbus_ARSIZE[2:0]),
       .dbus_ARBURST                    (dbus_ARBURST[1:0]),
       .dbus_ARLOCK                     (dbus_ARLOCK),
       .dbus_ARCACHE                    (dbus_ARCACHE[3:0]),
       .dbus_ARQOS                      (dbus_ARQOS[3:0]),
       .dbus_ARREGION                   (dbus_ARREGION[3:0]),
       .dbus_RREADY                     (dbus_RREADY),
       .dbus_AWVALID                    (dbus_AWVALID),
       .dbus_AWADDR                     (dbus_AWADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_AWPROT                     (dbus_AWPROT[2:0]),
       .dbus_AWID                       (dbus_AWID[AXI_ID_WIDTH-1:0]),
       .dbus_AWUSER                     (dbus_AWUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWLEN                      (dbus_AWLEN[7:0]),
       .dbus_AWSIZE                     (dbus_AWSIZE[2:0]),
       .dbus_AWBURST                    (dbus_AWBURST[1:0]),
       .dbus_AWLOCK                     (dbus_AWLOCK),
       .dbus_AWCACHE                    (dbus_AWCACHE[3:0]),
       .dbus_AWQOS                      (dbus_AWQOS[3:0]),
       .dbus_AWREGION                   (dbus_AWREGION[3:0]),
       .dbus_WVALID                     (dbus_WVALID),
       .dbus_WDATA                      (dbus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_WSTRB                      (dbus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]),
       .dbus_WLAST                      (dbus_WLAST),
       .dbus_WUSER                      (dbus_WUSER[AXI_USER_WIDTH-1:0]),
       .dbus_BREADY                     (dbus_BREADY),
       .clk                             (clk),
       .rst                             (rst),
       .ex_valid                        (ex_valid[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_alu_opc_bus                  (ex_alu_opc_bus[9 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_lpu_opc_bus                  (ex_lpu_opc_bus[5 *(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_epu_opc_bus                  (ex_epu_opc_bus[8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_bru_opc_bus                  (ex_bru_opc_bus[8*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_lsu_opc_bus                  (ex_lsu_opc_bus[7*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_bpu_upd                      (ex_bpu_upd[(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_pc                           (ex_pc[(CONFIG_AW-2 )*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_imm                          (ex_imm[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_operand1                     (ex_operand1[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_operand2                     (ex_operand2[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_rf_waddr                     (ex_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .ex_rf_we                        (ex_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .irqs                            (irqs[CONFIG_NUM_IRQ-1:0]),
       .msr_immid                       (msr_immid[CONFIG_DW-1:0]),
       .msr_icid                        (msr_icid[CONFIG_DW-1:0]),
       .msr_icinv_ready                 (msr_icinv_ready),
       .dbus_ARREADY                    (dbus_ARREADY),
       .dbus_RVALID                     (dbus_RVALID),
       .dbus_RDATA                      (dbus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_RRESP                      (dbus_RRESP[1:0]),
       .dbus_RLAST                      (dbus_RLAST),
       .dbus_RID                        (dbus_RID[AXI_ID_WIDTH-1:0]),
       .dbus_RUSER                      (dbus_RUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWREADY                    (dbus_AWREADY),
       .dbus_WREADY                     (dbus_WREADY),
       .dbus_BVALID                     (dbus_BVALID),
       .dbus_BRESP                      (dbus_BRESP[1:0]),
       .dbus_BID                        (dbus_BID[AXI_ID_WIDTH-1:0]),
       .dbus_BUSER                      (dbus_BUSER[AXI_USER_WIDTH-1:0]));
   ysyx_20210479_cmt
      #(
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH))
   U_CMT
      (
       .arf_RDATA                       (arf_RDATA[(1<<CONFIG_P_ISSUE_WIDTH)*2*CONFIG_DW-1:0]),
       .clk                             (clk),
       .commit_rf_wdat                  (commit_rf_wdat[CONFIG_DW*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .commit_rf_waddr                 (commit_rf_waddr[5*(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .commit_rf_we                    (commit_rf_we[(1<<CONFIG_P_ISSUE_WIDTH)-1:0]),
       .arf_RE                          (arf_RE[(1<<CONFIG_P_ISSUE_WIDTH)*2-1:0]),
       .arf_RADDR                       (arf_RADDR[(1<<CONFIG_P_ISSUE_WIDTH)*2*5-1:0]));
endmodule
module ysyx_20210479_prefetch_buf
#(
   parameter                           CONFIG_AW = 32,
   parameter                           CONFIG_P_FETCH_WIDTH = 2,
   parameter                           CONFIG_P_ISSUE_WIDTH = 2,
   parameter                           CONFIG_P_IQ_DEPTH = 4, 
   parameter                           CONFIG_PHT_P_NUM = 0,
   parameter                           CONFIG_BTB_P_NUM = 0
)
(
   input                               clk,
   input                               rst,
   input                               flush,
   input [((2 <<1)*8) * (1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_ins,
   input [(CONFIG_AW-2 ) * (1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_pc,
   input [2 * (1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_exc,
   input [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) * (1<<CONFIG_P_FETCH_WIDTH)-1:0] iq_bpu_upd,
   input [CONFIG_P_FETCH_WIDTH:0]      iq_push_cnt,
   input [CONFIG_P_FETCH_WIDTH:0]      iq_push_offset,
   output                              iq_ready,
   output [(1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_valid,
   input [CONFIG_P_ISSUE_WIDTH:0]      id_pop_cnt,
   output [((2 <<1)*8) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_ins,
   output [(CONFIG_AW-2 ) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_pc,
   output [2 * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_exc,
   output [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) * (1<<CONFIG_P_ISSUE_WIDTH)-1:0] id_bpu_upd
);
   localparam FW                       = (1<<CONFIG_P_FETCH_WIDTH);
   localparam IW                       = (1<<CONFIG_P_ISSUE_WIDTH);
   localparam FIFO_DW                  = (((2 <<1)*8) + (CONFIG_AW-2 ) + 2 + (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)); 
   localparam P_BANKS                  = (CONFIG_P_FETCH_WIDTH);
   localparam BANKS                    = (1<<P_BANKS);
   wire [P_BANKS-1:0]                  head_ff, tail_ff;
   wire [P_BANKS-1:0]                  head_nxt, tail_nxt;
   wire [P_BANKS-1:0]                  head_l                        [FW-1:0];
   wire [P_BANKS-1:0]                  head_r                        [FW-1:0];
   wire [P_BANKS-1:0]                  tail_r                        [FW-1:0];
   wire [P_BANKS-1:0]                  tail_inv                      [FW-1:0];
   wire [FIFO_DW-1:0]                  que_din                       [BANKS-1:0];
   wire [FIFO_DW-1:0]                  que_dout                      [BANKS-1:0];
   wire                                que_valid                     [BANKS-1:0];
   wire [BANKS-1:0]                    que_ready;
   wire                                que_push                      [BANKS-1:0];
   wire                                que_pop                       [BANKS-1:0];
   wire [((2 <<1)*8)-1:0]            iq_ins_unpacked               [FW-1:0];
   wire [(CONFIG_AW-2 )-1:0]                    iq_pc_unpacked                [FW-1:0];
   wire [2-1:0]               iq_exc_unpacked               [FW-1:0];
   wire [(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)-1:0]               iq_bpu_upd_unpacked           [FW-1:0];
   wire [P_BANKS:0]                    pop_cnt_adapt;
   genvar i;
   generate
      for(i=0;i<BANKS;i=i+1)
         begin : gen_ptr
            assign head_l[i]  = i + head_ff;
            assign head_r[i]  = i - head_ff;
            assign tail_r[i] = i - tail_ff;
            assign tail_inv[i] = i - tail_ff + iq_push_offset[P_BANKS-1:0];
         end
   endgenerate
   generate
      for(i=0;i<FW;i=i+1)
         begin
            assign iq_ins_unpacked[i] = iq_ins[i*((2 <<1)*8) +: ((2 <<1)*8)];
            assign iq_pc_unpacked[i] = iq_pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )];
            assign iq_exc_unpacked[i] = iq_exc[i*2 +: 2];
            assign iq_bpu_upd_unpacked[i] = iq_bpu_upd[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)];
         end
   endgenerate
   generate
      if (P_BANKS == CONFIG_P_ISSUE_WIDTH)
         assign pop_cnt_adapt = id_pop_cnt;
      else
         assign pop_cnt_adapt = {{P_BANKS-CONFIG_P_ISSUE_WIDTH{1'b0}}, id_pop_cnt};
   endgenerate
   generate
      for(i=0;i<BANKS;i=i+1)
         begin : gen_bank_ctrl
            assign que_din[i] = {iq_ins_unpacked[tail_inv[i]],
                                 iq_pc_unpacked[tail_inv[i]],
                                 iq_exc_unpacked[tail_inv[i]],
                                 iq_bpu_upd_unpacked[tail_inv[i]]};
            assign que_pop[i]  = ({1'b0, head_r[i]} < pop_cnt_adapt);
            assign que_push[i] = ({1'b0, tail_r[i]} < iq_push_cnt);
         end
   endgenerate
   assign head_nxt = (head_ff + pop_cnt_adapt[P_BANKS-1:0]) & {P_BANKS{~flush}};
   assign tail_nxt = (tail_ff + iq_push_cnt[P_BANKS-1:0]) & {P_BANKS{~flush}};
   ysyx_20210479_mDFF_r #(.DW(P_BANKS)) ff_head (.CLK(clk), .RST(rst), .D(head_nxt), .Q(head_ff) );
   ysyx_20210479_mDFF_r #(.DW(P_BANKS)) ff_tail (.CLK(clk), .RST(rst), .D(tail_nxt), .Q(tail_ff) );
   generate
      for(i=0;i<BANKS;i=i+1)
         begin
            ysyx_20210479_fifo_fwft
               #(
                  .DW            (FIFO_DW),
                  .DEPTH_WIDTH   (CONFIG_P_IQ_DEPTH)
               )
            U_FIFO
               (
                  .clk           (clk),
                  .rst           (rst),
                  .flush         (flush),
                  .push          (que_push[i]),
                  .din           (que_din[i]),
                  .ready         (que_ready[i]),
                  .pop           (que_pop[i]),
                  .dout          (que_dout[i]),
                  .valid         (que_valid[i])
               );
         end
   endgenerate
   generate
      for(i=0;i<(1<<CONFIG_P_ISSUE_WIDTH);i=i+1)
         begin : gen_pop
            assign {id_ins[i*((2 <<1)*8) +: ((2 <<1)*8)],
                     id_pc[i*(CONFIG_AW-2 ) +: (CONFIG_AW-2 )],
                     id_exc[i*2 +: 2],
                     id_bpu_upd[i*(2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1) +: (2 + CONFIG_PHT_P_NUM + CONFIG_BTB_P_NUM + (CONFIG_AW-2 ) + 1)] } = que_dout[head_l[i]];
            assign id_valid[i] = que_valid[head_l[i]];
         end
   endgenerate
   assign iq_ready = &que_ready;
endmodule
module ysyx_20210479_align_r
#(
   parameter                           AXI_P_DW_BYTES = 0,
   parameter                           PAYLOAD_P_DW_BYTES = 0,
   parameter                           RAM_AW = 0
)
(
   input [(1<<AXI_P_DW_BYTES)*8-1:0]   i_axi_RDATA,
   input                               i_ram_we,
   input [RAM_AW-1:0]                  i_ram_addr,
   output [(1<<PAYLOAD_P_DW_BYTES)-1:0] o_ram_wmsk,
   output [(1<<PAYLOAD_P_DW_BYTES)*8-1:0] o_ram_din
);
   localparam AXI_BYTES                = (1<<AXI_P_DW_BYTES);
   localparam PAYLOAD_BYTES            = (1<<PAYLOAD_P_DW_BYTES);
   genvar i;
   generate
      if (PAYLOAD_P_DW_BYTES == AXI_P_DW_BYTES)
         begin
            assign o_ram_din = i_axi_RDATA;
            assign o_ram_wmsk = {(1<<PAYLOAD_P_DW_BYTES){i_ram_we}};
         end
      else if (PAYLOAD_P_DW_BYTES < AXI_P_DW_BYTES)
         begin
            localparam WIN_NUM = (AXI_BYTES/PAYLOAD_BYTES);
            localparam WIN_P_NUM = (AXI_P_DW_BYTES - PAYLOAD_P_DW_BYTES);
            localparam WIN_DW = (PAYLOAD_BYTES*8);
            localparam WIN_P_DW_BYTES = (PAYLOAD_P_DW_BYTES);
            wire [WIN_DW-1:0] RDATA_win [WIN_NUM-1:0];
            for(i=0;i<WIN_NUM;i=i+1)
               assign RDATA_win[i] = i_axi_RDATA[i*WIN_DW +: WIN_DW];
            assign o_ram_din = RDATA_win[i_ram_addr[WIN_P_DW_BYTES +: WIN_P_NUM]];
            assign o_ram_wmsk = {(1<<PAYLOAD_P_DW_BYTES){i_ram_we}};
         end
      else
         begin
            localparam WIN_NUM = (PAYLOAD_BYTES/AXI_BYTES);
            localparam WIN_P_NUM = (PAYLOAD_P_DW_BYTES - AXI_P_DW_BYTES);
            localparam WIN_DW = (AXI_BYTES*8);
            localparam WIN_P_DW_BYTES = (AXI_P_DW_BYTES);
            wire [(1<<PAYLOAD_P_DW_BYTES)-1:0] ram_wmsk_tmp;
            for(i=0;i<WIN_NUM;i=i+1)
               assign ram_wmsk_tmp[i*(WIN_DW/8) +: (WIN_DW/8)] = {(WIN_DW/8){i_ram_addr[WIN_P_DW_BYTES +: WIN_P_NUM] == i}};
            assign o_ram_wmsk = ({(1<<PAYLOAD_P_DW_BYTES){i_ram_we}} & ram_wmsk_tmp);
            for(i=0;i<WIN_NUM;i=i+1)
               assign o_ram_din[i*WIN_DW +: WIN_DW] = i_axi_RDATA;
         end
   endgenerate
endmodule
module ysyx_20210479_align_w
#(
   parameter                           AXI_P_DW_BYTES = 0,
   parameter                           PAYLOAD_P_DW_BYTES = 0,
   parameter                           I_AXI_ADDR_AW = 0
)
(
   input [(1<<PAYLOAD_P_DW_BYTES)*8-1:0] i_axi_din,
   input                               i_axi_we,
   input [I_AXI_ADDR_AW-1:0]           i_axi_addr,
   output [(1<<AXI_P_DW_BYTES)-1:0]    o_axi_WSTRB,
   output [(1<<AXI_P_DW_BYTES)*8-1:0]  o_axi_WDATA
);
   localparam AXI_BYTES                = (1<<AXI_P_DW_BYTES);
   localparam PAYLOAD_BYTES            = (1<<PAYLOAD_P_DW_BYTES);
   genvar i;
   generate
      if (PAYLOAD_P_DW_BYTES == AXI_P_DW_BYTES)
         begin
            assign o_axi_WSTRB = {(1<<AXI_P_DW_BYTES){i_axi_we}};
            assign o_axi_WDATA = i_axi_din;
         end
      else if (PAYLOAD_P_DW_BYTES <= AXI_P_DW_BYTES)
         begin
            localparam WIN_NUM = (AXI_BYTES/PAYLOAD_BYTES);
            localparam WIN_P_NUM = (AXI_P_DW_BYTES - PAYLOAD_P_DW_BYTES);
            localparam WIN_DW = (PAYLOAD_BYTES*8);
            localparam WIN_P_DW_BYTES = (PAYLOAD_P_DW_BYTES);
            wire [(1<<AXI_P_DW_BYTES)-1:0] wstrb_tmp;
            for(i=0;i<WIN_NUM;i=i+1)
               assign wstrb_tmp[i*(WIN_DW/8) +: (WIN_DW/8)] = {(WIN_DW/8){i_axi_addr[WIN_P_DW_BYTES +: WIN_P_NUM] == i}};
            assign o_axi_WSTRB = ({(1<<AXI_P_DW_BYTES){i_axi_we}} & wstrb_tmp);
            for(i=0;i<WIN_NUM;i=i+1)
               assign o_axi_WDATA[i*WIN_DW +: WIN_DW] = i_axi_din;
         end
      else
         begin
            localparam WIN_NUM = (PAYLOAD_BYTES/AXI_BYTES);
            localparam WIN_P_NUM = (PAYLOAD_P_DW_BYTES - AXI_P_DW_BYTES);
            localparam WIN_DW = (AXI_BYTES*8);
            localparam WIN_P_DW_BYTES = (AXI_P_DW_BYTES);
            wire [WIN_DW-1:0] i_axi_din_win [WIN_NUM-1:0];
            for(i=0;i<WIN_NUM;i=i+1)
               assign i_axi_din_win[i] = i_axi_din[i*WIN_DW +: WIN_DW];
            assign o_axi_WDATA = i_axi_din_win[i_axi_addr[WIN_P_DW_BYTES +: WIN_P_NUM]];
            assign o_axi_WSTRB = {(1<<AXI_P_DW_BYTES){i_axi_we}};
         end
   endgenerate
endmodule
module ysyx_20210479_fifo_fwft
#(
   parameter DW = 8, 
   parameter DEPTH_WIDTH = 4 
)
(
   input                               clk,
   input                               rst,
   input                               flush,
   input                               push,
   input [DW-1:0]                      din,
   output                              ready,
   input                               pop,
   output [DW-1:0]                     dout,
   output                              valid
);
   wire [DEPTH_WIDTH:0]                ff_w_ptr;
   wire [DEPTH_WIDTH:0]                w_ptr_nxt;
   wire [DEPTH_WIDTH:0]                ff_r_ptr;
   wire [DEPTH_WIDTH:0]                r_ptr_nxt;
   wire [DW-1:0]                       rf_dout, rf_dout_byp;
   wire                                state_r;
   wire                                fwft_nxt;
   wire                                clr_state;
   wire [DW-1:0]                       dat_r, din_r;
   wire                                rf_conflict;
   wire                                rf_bypass;
   assign w_ptr_nxt = (ff_w_ptr + 1'd1) & {DEPTH_WIDTH+1{~flush}};
   assign r_ptr_nxt = (ff_r_ptr + 1'd1) & {DEPTH_WIDTH+1{~flush}};
   ysyx_20210479_mDFF_lr #(.DW(DEPTH_WIDTH + 1)) ff_w_ptr_r (.CLK(clk), .RST(rst), .LOAD(push|flush), .D(w_ptr_nxt), .Q(ff_w_ptr) );
   ysyx_20210479_mDFF_lr #(.DW(DEPTH_WIDTH + 1)) ff_r_ptr_r (.CLK(clk), .RST(rst), .LOAD(pop|flush), .D(r_ptr_nxt), .Q(ff_r_ptr) );
   assign ready = (ff_w_ptr[DEPTH_WIDTH] == ff_r_ptr[DEPTH_WIDTH]) |
                  (ff_w_ptr[DEPTH_WIDTH-1:0] != ff_r_ptr[DEPTH_WIDTH-1:0]); 
   assign valid = (ff_w_ptr != ff_r_ptr); 
   assign fwft_nxt = (~state_r & ~valid & push);
   assign clr_state = (state_r & pop);
   ysyx_20210479_mDFF_lr #(.DW(DW)) ff_dat (.CLK(clk), .RST(rst), .LOAD(fwft_nxt), .D(din), .Q(dat_r) );
   ysyx_20210479_mDFF_l #(.DW(DW)) ff_din (.CLK(clk), .LOAD(pop), .D(din), .Q(din_r) );
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_state (.CLK(clk),.RST(rst), .LOAD(fwft_nxt|clr_state|flush), .D((fwft_nxt|~clr_state) & ~flush), .Q(state_r) );
   assign dout = state_r ? dat_r : rf_dout_byp;
   ysyx_20210479_mRF_nwnr
      #(
         .DW (DW),
         .AW (DEPTH_WIDTH),
         .NUM_READ   (1),
         .NUM_WRITE  (1)
      )
   U_RF
      (
         .CLK     (clk),
         .RE      (pop),
         .RADDR   (r_ptr_nxt[DEPTH_WIDTH-1:0]),
         .RDATA   (rf_dout),
         .WE      (push),
         .WADDR   (ff_w_ptr[DEPTH_WIDTH-1:0]),
         .WDATA   (din)
      );
   assign rf_conflict = ((ff_w_ptr[DEPTH_WIDTH-1:0] == r_ptr_nxt[DEPTH_WIDTH-1:0]) & push & pop);
   ysyx_20210479_mDFF_lr #(.DW(1)) ff_bypass (.CLK(clk), .RST(rst), .LOAD(rf_conflict | pop), .D(rf_conflict | ~pop), .Q(rf_bypass) );
   assign rf_dout_byp = rf_bypass ? din_r : rf_dout;
endmodule
module ysyx_20210479_pmux
#(
   parameter SELW = 0,
   parameter DW = 0
)
(
   input [SELW-1:0] sel,
   input [DW*SELW-1:0] din,
   output reg [DW-1:0] dout
);
   generate
      if (SELW==2)
         begin : gen_enc_2
            always @(*)
                begin
                    casez(sel)
                       2'b?1: dout = din[0*DW +: DW];
                       2'b10: dout = din[1*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==3)
         begin : gen_enc_3
            always @(*)
                begin
                    casez(sel)
                       3'b??1: dout = din[0*DW +: DW];
                       3'b?10: dout = din[1*DW +: DW];
                       3'b100: dout = din[2*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==4)
         begin : gen_enc_4
            always @(*)
                begin
                    casez(sel)
                       4'b???1: dout = din[0*DW +: DW];
                       4'b??10: dout = din[1*DW +: DW];
                       4'b?100: dout = din[2*DW +: DW];
                       4'b1000: dout = din[3*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==5)
         begin : gen_enc_5
            always @(*)
                begin
                    casez(sel)
                       5'b????1: dout = din[0*DW +: DW];
                       5'b???10: dout = din[1*DW +: DW];
                       5'b??100: dout = din[2*DW +: DW];
                       5'b?1000: dout = din[3*DW +: DW];
                       5'b10000: dout = din[4*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==6)
         begin : gen_enc_6
            always @(*)
                begin
                    casez(sel)
                       6'b?????1: dout = din[0*DW +: DW];
                       6'b????10: dout = din[1*DW +: DW];
                       6'b???100: dout = din[2*DW +: DW];
                       6'b??1000: dout = din[3*DW +: DW];
                       6'b?10000: dout = din[4*DW +: DW];
                       6'b100000: dout = din[5*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==7)
         begin : gen_enc_7
            always @(*)
                begin
                    casez(sel)
                       7'b??????1: dout = din[0*DW +: DW];
                       7'b?????10: dout = din[1*DW +: DW];
                       7'b????100: dout = din[2*DW +: DW];
                       7'b???1000: dout = din[3*DW +: DW];
                       7'b??10000: dout = din[4*DW +: DW];
                       7'b?100000: dout = din[5*DW +: DW];
                       7'b1000000: dout = din[6*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==8)
         begin : gen_enc_8
            always @(*)
                begin
                    casez(sel)
                       8'b???????1: dout = din[0*DW +: DW];
                       8'b??????10: dout = din[1*DW +: DW];
                       8'b?????100: dout = din[2*DW +: DW];
                       8'b????1000: dout = din[3*DW +: DW];
                       8'b???10000: dout = din[4*DW +: DW];
                       8'b??100000: dout = din[5*DW +: DW];
                       8'b?1000000: dout = din[6*DW +: DW];
                       8'b10000000: dout = din[7*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      if (SELW==9)
         begin : gen_enc_9
            always @(*)
                begin
                    casez(sel)
                       9'b????????1: dout = din[0*DW +: DW];
                       9'b???????10: dout = din[1*DW +: DW];
                       9'b??????100: dout = din[2*DW +: DW];
                       9'b?????1000: dout = din[3*DW +: DW];
                       9'b????10000: dout = din[4*DW +: DW];
                       9'b???100000: dout = din[5*DW +: DW];
                       9'b??1000000: dout = din[6*DW +: DW];
                       9'b?10000000: dout = din[7*DW +: DW];
                       9'b100000000: dout = din[8*DW +: DW];
                       default: begin dout = din[0 +: DW]; end
                    endcase
                end
         end
      else
      begin : gen_enc_fail
            initial
                $fatal("\n Unimplemented size. Please update parameters of generator. \n");
         end
    endgenerate
endmodule
module ysyx_20210479_pmux_v
#(
   parameter SELW = 0,
   parameter DW = 0
)
(
   input [SELW-1:0] sel,
   input [DW*SELW-1:0] din,
   output reg [DW-1:0] dout
   , output reg valid
);
   generate
      if (SELW==2)
         begin : gen_enc_2
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       2'b?1: dout = din[0*DW +: DW];
                       2'b10: dout = din[1*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==3)
         begin : gen_enc_3
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       3'b??1: dout = din[0*DW +: DW];
                       3'b?10: dout = din[1*DW +: DW];
                       3'b100: dout = din[2*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==4)
         begin : gen_enc_4
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       4'b???1: dout = din[0*DW +: DW];
                       4'b??10: dout = din[1*DW +: DW];
                       4'b?100: dout = din[2*DW +: DW];
                       4'b1000: dout = din[3*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==5)
         begin : gen_enc_5
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       5'b????1: dout = din[0*DW +: DW];
                       5'b???10: dout = din[1*DW +: DW];
                       5'b??100: dout = din[2*DW +: DW];
                       5'b?1000: dout = din[3*DW +: DW];
                       5'b10000: dout = din[4*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==6)
         begin : gen_enc_6
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       6'b?????1: dout = din[0*DW +: DW];
                       6'b????10: dout = din[1*DW +: DW];
                       6'b???100: dout = din[2*DW +: DW];
                       6'b??1000: dout = din[3*DW +: DW];
                       6'b?10000: dout = din[4*DW +: DW];
                       6'b100000: dout = din[5*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==7)
         begin : gen_enc_7
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       7'b??????1: dout = din[0*DW +: DW];
                       7'b?????10: dout = din[1*DW +: DW];
                       7'b????100: dout = din[2*DW +: DW];
                       7'b???1000: dout = din[3*DW +: DW];
                       7'b??10000: dout = din[4*DW +: DW];
                       7'b?100000: dout = din[5*DW +: DW];
                       7'b1000000: dout = din[6*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==8)
         begin : gen_enc_8
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       8'b???????1: dout = din[0*DW +: DW];
                       8'b??????10: dout = din[1*DW +: DW];
                       8'b?????100: dout = din[2*DW +: DW];
                       8'b????1000: dout = din[3*DW +: DW];
                       8'b???10000: dout = din[4*DW +: DW];
                       8'b??100000: dout = din[5*DW +: DW];
                       8'b?1000000: dout = din[6*DW +: DW];
                       8'b10000000: dout = din[7*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      if (SELW==9)
         begin : gen_enc_9
            always @(*)
                begin
                    valid = 'b1;
                    casez(sel)
                       9'b????????1: dout = din[0*DW +: DW];
                       9'b???????10: dout = din[1*DW +: DW];
                       9'b??????100: dout = din[2*DW +: DW];
                       9'b?????1000: dout = din[3*DW +: DW];
                       9'b????10000: dout = din[4*DW +: DW];
                       9'b???100000: dout = din[5*DW +: DW];
                       9'b??1000000: dout = din[6*DW +: DW];
                       9'b?10000000: dout = din[7*DW +: DW];
                       9'b100000000: dout = din[8*DW +: DW];
                       default: begin dout = din[0 +: DW]; valid = 'b0; end
                    endcase
                end
         end
      else
      begin : gen_enc_fail
            initial
                $fatal("\n Unimplemented size. Please update parameters of generator. \n");
         end
    endgenerate
endmodule
module ysyx_20210479_popcnt
#(
   parameter DW = 0,
   parameter P_DW = 0 
)
(
   input [DW-1:0] bitmap,
   output reg [P_DW:0] count
);
   integer j;
   always @(*)
      begin
         count = 'b0;
         for(j=0;j<(1<<P_DW);j=j+1)
            count = count + {{P_DW{1'b0}}, bitmap[j]};
      end
endmodule
module ysyx_20210479_priority_encoder
#(
   parameter P_DW = 0
)
(
   input [(1<<P_DW)-1:0] din,
   output reg [P_DW-1:0] dout
);
   generate
      if (P_DW==1)
        begin : gen_enc_1
            always @(*)
                begin
                    casez(din)
                       2'b?1: dout = 1'd0;
                       2'b10: dout = 1'd1;
                       default: begin dout = 1'd0; end
                    endcase
                end
        end
      else if (P_DW==2)
        begin : gen_enc_2
            always @(*)
                begin
                    casez(din)
                       4'b???1: dout = 2'd0;
                       4'b??10: dout = 2'd1;
                       4'b?100: dout = 2'd2;
                       4'b1000: dout = 2'd3;
                       default: begin dout = 2'd0; end
                    endcase
                end
        end
      else if (P_DW==3)
        begin : gen_enc_3
            always @(*)
                begin
                    casez(din)
                       8'b???????1: dout = 3'd0;
                       8'b??????10: dout = 3'd1;
                       8'b?????100: dout = 3'd2;
                       8'b????1000: dout = 3'd3;
                       8'b???10000: dout = 3'd4;
                       8'b??100000: dout = 3'd5;
                       8'b?1000000: dout = 3'd6;
                       8'b10000000: dout = 3'd7;
                       default: begin dout = 3'd0; end
                    endcase
                end
        end
      else if (P_DW==4)
        begin : gen_enc_4
            always @(*)
                begin
                    casez(din)
                       16'b???????????????1: dout = 4'd0;
                       16'b??????????????10: dout = 4'd1;
                       16'b?????????????100: dout = 4'd2;
                       16'b????????????1000: dout = 4'd3;
                       16'b???????????10000: dout = 4'd4;
                       16'b??????????100000: dout = 4'd5;
                       16'b?????????1000000: dout = 4'd6;
                       16'b????????10000000: dout = 4'd7;
                       16'b???????100000000: dout = 4'd8;
                       16'b??????1000000000: dout = 4'd9;
                       16'b?????10000000000: dout = 4'd10;
                       16'b????100000000000: dout = 4'd11;
                       16'b???1000000000000: dout = 4'd12;
                       16'b??10000000000000: dout = 4'd13;
                       16'b?100000000000000: dout = 4'd14;
                       16'b1000000000000000: dout = 4'd15;
                       default: begin dout = 4'd0; end
                    endcase
                end
        end
      else if (P_DW==5)
        begin : gen_enc_5
            always @(*)
                begin
                    casez(din)
                       32'b???????????????????????????????1: dout = 5'd0;
                       32'b??????????????????????????????10: dout = 5'd1;
                       32'b?????????????????????????????100: dout = 5'd2;
                       32'b????????????????????????????1000: dout = 5'd3;
                       32'b???????????????????????????10000: dout = 5'd4;
                       32'b??????????????????????????100000: dout = 5'd5;
                       32'b?????????????????????????1000000: dout = 5'd6;
                       32'b????????????????????????10000000: dout = 5'd7;
                       32'b???????????????????????100000000: dout = 5'd8;
                       32'b??????????????????????1000000000: dout = 5'd9;
                       32'b?????????????????????10000000000: dout = 5'd10;
                       32'b????????????????????100000000000: dout = 5'd11;
                       32'b???????????????????1000000000000: dout = 5'd12;
                       32'b??????????????????10000000000000: dout = 5'd13;
                       32'b?????????????????100000000000000: dout = 5'd14;
                       32'b????????????????1000000000000000: dout = 5'd15;
                       32'b???????????????10000000000000000: dout = 5'd16;
                       32'b??????????????100000000000000000: dout = 5'd17;
                       32'b?????????????1000000000000000000: dout = 5'd18;
                       32'b????????????10000000000000000000: dout = 5'd19;
                       32'b???????????100000000000000000000: dout = 5'd20;
                       32'b??????????1000000000000000000000: dout = 5'd21;
                       32'b?????????10000000000000000000000: dout = 5'd22;
                       32'b????????100000000000000000000000: dout = 5'd23;
                       32'b???????1000000000000000000000000: dout = 5'd24;
                       32'b??????10000000000000000000000000: dout = 5'd25;
                       32'b?????100000000000000000000000000: dout = 5'd26;
                       32'b????1000000000000000000000000000: dout = 5'd27;
                       32'b???10000000000000000000000000000: dout = 5'd28;
                       32'b??100000000000000000000000000000: dout = 5'd29;
                       32'b?1000000000000000000000000000000: dout = 5'd30;
                       32'b10000000000000000000000000000000: dout = 5'd31;
                       default: begin dout = 5'd0; end
                    endcase
                end
        end
      else if (P_DW==6)
        begin : gen_enc_6
            always @(*)
                begin
                    casez(din)
                       64'b???????????????????????????????????????????????????????????????1: dout = 6'd0;
                       64'b??????????????????????????????????????????????????????????????10: dout = 6'd1;
                       64'b?????????????????????????????????????????????????????????????100: dout = 6'd2;
                       64'b????????????????????????????????????????????????????????????1000: dout = 6'd3;
                       64'b???????????????????????????????????????????????????????????10000: dout = 6'd4;
                       64'b??????????????????????????????????????????????????????????100000: dout = 6'd5;
                       64'b?????????????????????????????????????????????????????????1000000: dout = 6'd6;
                       64'b????????????????????????????????????????????????????????10000000: dout = 6'd7;
                       64'b???????????????????????????????????????????????????????100000000: dout = 6'd8;
                       64'b??????????????????????????????????????????????????????1000000000: dout = 6'd9;
                       64'b?????????????????????????????????????????????????????10000000000: dout = 6'd10;
                       64'b????????????????????????????????????????????????????100000000000: dout = 6'd11;
                       64'b???????????????????????????????????????????????????1000000000000: dout = 6'd12;
                       64'b??????????????????????????????????????????????????10000000000000: dout = 6'd13;
                       64'b?????????????????????????????????????????????????100000000000000: dout = 6'd14;
                       64'b????????????????????????????????????????????????1000000000000000: dout = 6'd15;
                       64'b???????????????????????????????????????????????10000000000000000: dout = 6'd16;
                       64'b??????????????????????????????????????????????100000000000000000: dout = 6'd17;
                       64'b?????????????????????????????????????????????1000000000000000000: dout = 6'd18;
                       64'b????????????????????????????????????????????10000000000000000000: dout = 6'd19;
                       64'b???????????????????????????????????????????100000000000000000000: dout = 6'd20;
                       64'b??????????????????????????????????????????1000000000000000000000: dout = 6'd21;
                       64'b?????????????????????????????????????????10000000000000000000000: dout = 6'd22;
                       64'b????????????????????????????????????????100000000000000000000000: dout = 6'd23;
                       64'b???????????????????????????????????????1000000000000000000000000: dout = 6'd24;
                       64'b??????????????????????????????????????10000000000000000000000000: dout = 6'd25;
                       64'b?????????????????????????????????????100000000000000000000000000: dout = 6'd26;
                       64'b????????????????????????????????????1000000000000000000000000000: dout = 6'd27;
                       64'b???????????????????????????????????10000000000000000000000000000: dout = 6'd28;
                       64'b??????????????????????????????????100000000000000000000000000000: dout = 6'd29;
                       64'b?????????????????????????????????1000000000000000000000000000000: dout = 6'd30;
                       64'b????????????????????????????????10000000000000000000000000000000: dout = 6'd31;
                       64'b???????????????????????????????100000000000000000000000000000000: dout = 6'd32;
                       64'b??????????????????????????????1000000000000000000000000000000000: dout = 6'd33;
                       64'b?????????????????????????????10000000000000000000000000000000000: dout = 6'd34;
                       64'b????????????????????????????100000000000000000000000000000000000: dout = 6'd35;
                       64'b???????????????????????????1000000000000000000000000000000000000: dout = 6'd36;
                       64'b??????????????????????????10000000000000000000000000000000000000: dout = 6'd37;
                       64'b?????????????????????????100000000000000000000000000000000000000: dout = 6'd38;
                       64'b????????????????????????1000000000000000000000000000000000000000: dout = 6'd39;
                       64'b???????????????????????10000000000000000000000000000000000000000: dout = 6'd40;
                       64'b??????????????????????100000000000000000000000000000000000000000: dout = 6'd41;
                       64'b?????????????????????1000000000000000000000000000000000000000000: dout = 6'd42;
                       64'b????????????????????10000000000000000000000000000000000000000000: dout = 6'd43;
                       64'b???????????????????100000000000000000000000000000000000000000000: dout = 6'd44;
                       64'b??????????????????1000000000000000000000000000000000000000000000: dout = 6'd45;
                       64'b?????????????????10000000000000000000000000000000000000000000000: dout = 6'd46;
                       64'b????????????????100000000000000000000000000000000000000000000000: dout = 6'd47;
                       64'b???????????????1000000000000000000000000000000000000000000000000: dout = 6'd48;
                       64'b??????????????10000000000000000000000000000000000000000000000000: dout = 6'd49;
                       64'b?????????????100000000000000000000000000000000000000000000000000: dout = 6'd50;
                       64'b????????????1000000000000000000000000000000000000000000000000000: dout = 6'd51;
                       64'b???????????10000000000000000000000000000000000000000000000000000: dout = 6'd52;
                       64'b??????????100000000000000000000000000000000000000000000000000000: dout = 6'd53;
                       64'b?????????1000000000000000000000000000000000000000000000000000000: dout = 6'd54;
                       64'b????????10000000000000000000000000000000000000000000000000000000: dout = 6'd55;
                       64'b???????100000000000000000000000000000000000000000000000000000000: dout = 6'd56;
                       64'b??????1000000000000000000000000000000000000000000000000000000000: dout = 6'd57;
                       64'b?????10000000000000000000000000000000000000000000000000000000000: dout = 6'd58;
                       64'b????100000000000000000000000000000000000000000000000000000000000: dout = 6'd59;
                       64'b???1000000000000000000000000000000000000000000000000000000000000: dout = 6'd60;
                       64'b??10000000000000000000000000000000000000000000000000000000000000: dout = 6'd61;
                       64'b?100000000000000000000000000000000000000000000000000000000000000: dout = 6'd62;
                       64'b1000000000000000000000000000000000000000000000000000000000000000: dout = 6'd63;
                       default: begin dout = 6'd0; end
                    endcase
                end
        end
      else if (P_DW==7)
        begin : gen_enc_7
            always @(*)
                begin
                    casez(din)
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1: dout = 7'd0;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10: dout = 7'd1;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100: dout = 7'd2;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000: dout = 7'd3;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000: dout = 7'd4;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000: dout = 7'd5;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000: dout = 7'd6;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000: dout = 7'd7;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000: dout = 7'd8;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000: dout = 7'd9;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000: dout = 7'd10;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000: dout = 7'd11;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000: dout = 7'd12;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000: dout = 7'd13;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000: dout = 7'd14;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000: dout = 7'd15;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000: dout = 7'd16;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000: dout = 7'd17;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000: dout = 7'd18;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000: dout = 7'd19;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000: dout = 7'd20;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000: dout = 7'd21;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000: dout = 7'd22;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000: dout = 7'd23;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000: dout = 7'd24;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000: dout = 7'd25;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000: dout = 7'd26;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000: dout = 7'd27;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000: dout = 7'd28;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000: dout = 7'd29;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000: dout = 7'd30;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000: dout = 7'd31;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000: dout = 7'd32;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000: dout = 7'd33;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000: dout = 7'd34;
                       128'b????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000: dout = 7'd35;
                       128'b???????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000: dout = 7'd36;
                       128'b??????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000: dout = 7'd37;
                       128'b?????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000: dout = 7'd38;
                       128'b????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000: dout = 7'd39;
                       128'b???????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000: dout = 7'd40;
                       128'b??????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000: dout = 7'd41;
                       128'b?????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000: dout = 7'd42;
                       128'b????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000: dout = 7'd43;
                       128'b???????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000: dout = 7'd44;
                       128'b??????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000: dout = 7'd45;
                       128'b?????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000: dout = 7'd46;
                       128'b????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000: dout = 7'd47;
                       128'b???????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000: dout = 7'd48;
                       128'b??????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000: dout = 7'd49;
                       128'b?????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000: dout = 7'd50;
                       128'b????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000: dout = 7'd51;
                       128'b???????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000: dout = 7'd52;
                       128'b??????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000: dout = 7'd53;
                       128'b?????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000: dout = 7'd54;
                       128'b????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000: dout = 7'd55;
                       128'b???????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000: dout = 7'd56;
                       128'b??????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000: dout = 7'd57;
                       128'b?????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000: dout = 7'd58;
                       128'b????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000: dout = 7'd59;
                       128'b???????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000: dout = 7'd60;
                       128'b??????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000: dout = 7'd61;
                       128'b?????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000: dout = 7'd62;
                       128'b????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000: dout = 7'd63;
                       128'b???????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000: dout = 7'd64;
                       128'b??????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000: dout = 7'd65;
                       128'b?????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd66;
                       128'b????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd67;
                       128'b???????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd68;
                       128'b??????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd69;
                       128'b?????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd70;
                       128'b????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd71;
                       128'b???????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd72;
                       128'b??????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd73;
                       128'b?????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd74;
                       128'b????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd75;
                       128'b???????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd76;
                       128'b??????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd77;
                       128'b?????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd78;
                       128'b????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd79;
                       128'b???????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd80;
                       128'b??????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd81;
                       128'b?????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd82;
                       128'b????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd83;
                       128'b???????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd84;
                       128'b??????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd85;
                       128'b?????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd86;
                       128'b????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd87;
                       128'b???????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd88;
                       128'b??????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd89;
                       128'b?????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd90;
                       128'b????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd91;
                       128'b???????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd92;
                       128'b??????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd93;
                       128'b?????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd94;
                       128'b????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd95;
                       128'b???????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd96;
                       128'b??????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd97;
                       128'b?????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd98;
                       128'b????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd99;
                       128'b???????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd100;
                       128'b??????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd101;
                       128'b?????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd102;
                       128'b????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd103;
                       128'b???????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd104;
                       128'b??????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd105;
                       128'b?????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd106;
                       128'b????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd107;
                       128'b???????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd108;
                       128'b??????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd109;
                       128'b?????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd110;
                       128'b????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd111;
                       128'b???????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd112;
                       128'b??????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd113;
                       128'b?????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd114;
                       128'b????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd115;
                       128'b???????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd116;
                       128'b??????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd117;
                       128'b?????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd118;
                       128'b????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd119;
                       128'b???????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd120;
                       128'b??????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd121;
                       128'b?????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd122;
                       128'b????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd123;
                       128'b???10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd124;
                       128'b??100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd125;
                       128'b?1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd126;
                       128'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 7'd127;
                       default: begin dout = 7'd0; end
                    endcase
                end
        end
      else if (P_DW==8)
        begin : gen_enc_8
            always @(*)
                begin
                    casez(din)
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1: dout = 8'd0;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10: dout = 8'd1;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100: dout = 8'd2;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000: dout = 8'd3;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000: dout = 8'd4;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000: dout = 8'd5;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000: dout = 8'd6;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000: dout = 8'd7;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000: dout = 8'd8;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000: dout = 8'd9;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000: dout = 8'd10;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000: dout = 8'd11;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000: dout = 8'd12;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000: dout = 8'd13;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000: dout = 8'd14;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000: dout = 8'd15;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000: dout = 8'd16;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000: dout = 8'd17;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000: dout = 8'd18;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000: dout = 8'd19;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000: dout = 8'd20;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000: dout = 8'd21;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000: dout = 8'd22;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000: dout = 8'd23;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000: dout = 8'd24;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000: dout = 8'd25;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000: dout = 8'd26;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000: dout = 8'd27;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000: dout = 8'd28;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000: dout = 8'd29;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000: dout = 8'd30;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000: dout = 8'd31;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000: dout = 8'd32;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000: dout = 8'd33;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000: dout = 8'd34;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000: dout = 8'd35;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000: dout = 8'd36;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000: dout = 8'd37;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000: dout = 8'd38;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000: dout = 8'd39;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000: dout = 8'd40;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000: dout = 8'd41;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000: dout = 8'd42;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000: dout = 8'd43;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000: dout = 8'd44;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000: dout = 8'd45;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000: dout = 8'd46;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000: dout = 8'd47;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000: dout = 8'd48;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000: dout = 8'd49;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000: dout = 8'd50;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000: dout = 8'd51;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000: dout = 8'd52;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000: dout = 8'd53;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000: dout = 8'd54;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000: dout = 8'd55;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000: dout = 8'd56;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000: dout = 8'd57;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000: dout = 8'd58;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000: dout = 8'd59;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000: dout = 8'd60;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000: dout = 8'd61;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000: dout = 8'd62;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000: dout = 8'd63;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000: dout = 8'd64;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000: dout = 8'd65;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd66;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd67;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd68;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd69;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd70;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd71;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd72;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd73;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd74;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd75;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd76;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd77;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd78;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd79;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd80;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd81;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd82;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd83;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd84;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd85;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd86;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd87;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd88;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd89;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd90;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd91;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd92;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd93;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd94;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd95;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd96;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd97;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd98;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd99;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd100;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd101;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd102;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd103;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd104;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd105;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd106;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd107;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd108;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd109;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd110;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd111;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd112;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd113;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd114;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd115;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd116;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd117;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd118;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd119;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd120;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd121;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd122;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd123;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd124;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd125;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd126;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd127;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd128;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd129;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd130;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd131;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd132;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd133;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd134;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd135;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd136;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd137;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd138;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd139;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd140;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd141;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd142;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd143;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd144;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd145;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd146;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd147;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd148;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd149;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd150;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd151;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd152;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd153;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd154;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd155;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd156;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd157;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd158;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd159;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd160;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd161;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd162;
                       256'b????????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd163;
                       256'b???????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd164;
                       256'b??????????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd165;
                       256'b?????????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd166;
                       256'b????????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd167;
                       256'b???????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd168;
                       256'b??????????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd169;
                       256'b?????????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd170;
                       256'b????????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd171;
                       256'b???????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd172;
                       256'b??????????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd173;
                       256'b?????????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd174;
                       256'b????????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd175;
                       256'b???????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd176;
                       256'b??????????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd177;
                       256'b?????????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd178;
                       256'b????????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd179;
                       256'b???????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd180;
                       256'b??????????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd181;
                       256'b?????????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd182;
                       256'b????????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd183;
                       256'b???????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd184;
                       256'b??????????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd185;
                       256'b?????????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd186;
                       256'b????????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd187;
                       256'b???????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd188;
                       256'b??????????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd189;
                       256'b?????????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd190;
                       256'b????????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd191;
                       256'b???????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd192;
                       256'b??????????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd193;
                       256'b?????????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd194;
                       256'b????????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd195;
                       256'b???????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd196;
                       256'b??????????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd197;
                       256'b?????????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd198;
                       256'b????????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd199;
                       256'b???????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd200;
                       256'b??????????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd201;
                       256'b?????????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd202;
                       256'b????????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd203;
                       256'b???????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd204;
                       256'b??????????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd205;
                       256'b?????????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd206;
                       256'b????????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd207;
                       256'b???????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd208;
                       256'b??????????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd209;
                       256'b?????????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd210;
                       256'b????????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd211;
                       256'b???????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd212;
                       256'b??????????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd213;
                       256'b?????????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd214;
                       256'b????????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd215;
                       256'b???????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd216;
                       256'b??????????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd217;
                       256'b?????????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd218;
                       256'b????????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd219;
                       256'b???????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd220;
                       256'b??????????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd221;
                       256'b?????????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd222;
                       256'b????????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd223;
                       256'b???????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd224;
                       256'b??????????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd225;
                       256'b?????????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd226;
                       256'b????????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd227;
                       256'b???????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd228;
                       256'b??????????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd229;
                       256'b?????????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd230;
                       256'b????????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd231;
                       256'b???????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd232;
                       256'b??????????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd233;
                       256'b?????????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd234;
                       256'b????????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd235;
                       256'b???????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd236;
                       256'b??????????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd237;
                       256'b?????????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd238;
                       256'b????????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd239;
                       256'b???????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd240;
                       256'b??????????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd241;
                       256'b?????????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd242;
                       256'b????????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd243;
                       256'b???????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd244;
                       256'b??????????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd245;
                       256'b?????????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd246;
                       256'b????????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd247;
                       256'b???????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd248;
                       256'b??????1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd249;
                       256'b?????10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd250;
                       256'b????100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd251;
                       256'b???1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd252;
                       256'b??10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd253;
                       256'b?100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd254;
                       256'b1000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000: dout = 8'd255;
                       default: begin dout = 8'd0; end
                    endcase
                end
        end
      else 
         begin : gen_enc_fail
            initial
                $fatal("\n Unimplemented size of binary encoder. Please update parameters of generator. \n");
         end
    endgenerate
endmodule
module ysyx_20210479_mDFF # (
   parameter DW = 1 
)
(
   input CLK,
   input [DW-1:0] D, 
   output reg [DW-1:0] Q 
);
   always @(posedge CLK)
      Q <= D;
endmodule
module ysyx_20210479_mDFF_l # (
   parameter DW = 1 
)
(
   input CLK,
   input LOAD,
   input [DW-1:0] D, 
   output reg [DW-1:0] Q 
);
   always @(posedge CLK)
      if (LOAD)
         Q <= D;
endmodule
module ysyx_20210479_mDFF_lr # (
   parameter DW = 1, 
   parameter RST_VECTOR = {DW{1'b0}}
)
(
   input CLK,
   input RST,
   input LOAD,
   input [DW-1:0] D, 
   output reg [DW-1:0] Q 
);
   always @(posedge CLK) begin
      if (RST)
         Q <= RST_VECTOR;
      else if (LOAD)
         Q <= D;
   end
endmodule
module ysyx_20210479_mDFF_r # (
   parameter DW = 1, 
   parameter RST_VECTOR = {DW{1'b0}}
)
(
   input CLK,
   input RST,
   input [DW-1:0] D, 
   output reg [DW-1:0] Q 
);
   always @(posedge CLK) begin
      if (RST)
         Q <= RST_VECTOR;
      else
         Q <= D;
   end
endmodule
module ysyx_20210479_mRAM_s_s_be
#(
   parameter P_DW = 0,
   parameter AW = 0
)
(
   input CLK,
   input [AW-1:0] ADDR,
   input RE,
   output [(1<<P_DW)-1:0] DOUT,
   input [(1<<P_DW)/8-1:0] WE,
   input [(1<<P_DW)-1:0] DIN
);
   localparam P_DW_BYTES = (P_DW-3);
   localparam SRAM_DW = 128;
   localparam SRAM_AW = 6;
   localparam SRAM_P_DW_BYTES = 4; 
   wire [(1<<P_DW)-1:0] we_bmsk;
   wire [AW-1:0] re_addr_ff;
   wire [AW-1:0] addr_w;
   genvar i;
   ysyx_20210479_mDFF_l #(.DW(AW)) ff_re_addr (.CLK(CLK), .LOAD(RE), .D(ADDR), .Q(re_addr_ff) );
   assign addr_w = (RE | (|WE)) ? ADDR : re_addr_ff;
   for(i=0;i<(1<<P_DW_BYTES);i=i+1)
      assign we_bmsk[i*8 +: 8] = {8{WE[i]}};
   generate
      if (((1<<P_DW) == SRAM_DW) && (AW == SRAM_AW))
         begin
            S011HD1P_X32Y2D128_BW U_S011HD1P_X32Y2D128_BW
               (
                  .Q                      (DOUT),
                  .CLK                    (CLK),
                  .CEN                    (1'b0),     
                  .WEN                    (~|WE),     
                  .BWEN                   (~we_bmsk), 
                  .A                      (addr_w),
                  .D                      (DIN)
               );
         end
      else if (((1<<P_DW) < SRAM_DW) && ((AW-(SRAM_P_DW_BYTES - P_DW_BYTES)) == SRAM_AW))
         begin
            localparam WIN_P_NUM = (SRAM_P_DW_BYTES - P_DW_BYTES);
            localparam WIN_NUM = (1<<WIN_P_NUM);
            localparam WIN_DW = (1<<P_DW);
            wire [SRAM_DW-1:0] sram_q;
            wire [SRAM_DW-1:0] sram_bwen;
            wire [SRAM_DW-1:0] sram_d;
            wire [WIN_DW-1:0] DOUT_win [WIN_NUM-1:0];
            for(i=0;i<WIN_NUM;i=i+1)
               assign sram_bwen[i*WIN_DW +: WIN_DW] = (we_bmsk & {WIN_DW{addr_w[WIN_P_NUM-1:0] == i}});
            for(i=0;i<WIN_NUM;i=i+1)
               assign sram_d[i*WIN_DW +: WIN_DW] = DIN;
            S011HD1P_X32Y2D128_BW S011HD1P_X32Y2D128_BW
               (
                  .Q                      (sram_q),
                  .CLK                    (CLK),
                  .CEN                    (1'b0),        
                  .WEN                    (~|WE),        
                  .BWEN                   (~sram_bwen),  
                  .A                      (addr_w[WIN_P_NUM +: SRAM_AW]),
                  .D                      (sram_d)
               );
            for(i=0;i<WIN_NUM;i=i+1)
               assign DOUT_win[i] = sram_q[i*WIN_DW +: WIN_DW];
            assign DOUT = DOUT_win[re_addr_ff[WIN_P_NUM-1:0]];
         end
      else
         begin
            initial $fatal(1, "SRAM with the specified size is unsupported.");
         end
   endgenerate
endmodule
module ysyx_20210479_mRF_1wr
#(
   parameter DW = 0,
   parameter AW = 0
)
(
   input CLK,
   input [AW-1:0] ADDR,
   input RE,
   output [DW-1:0] RDATA,
   input WE,
   input [DW-1:0] WDATA
);
   reg [DW-1:0] regfile [(1<<AW)-1:0];
   reg [DW-1:0] ff_dout;
   always @(posedge CLK)
      begin
         if (WE)
            regfile[ADDR] <= WDATA;
         if (RE)
            ff_dout <= regfile[ADDR];
      end
   assign RDATA = ff_dout;
endmodule
module ysyx_20210479_mRF_nwnr
#(
   parameter DW = 0,
   parameter AW = 0,
   parameter NUM_READ = 0,
   parameter NUM_WRITE = 0
)
(
   input CLK,
   input [NUM_READ-1:0] RE,
   input [NUM_READ*AW-1:0] RADDR,
   output [NUM_READ*DW-1:0] RDATA,
   input [NUM_WRITE-1:0] WE,
   input [AW*NUM_WRITE-1:0] WADDR,
   input [DW*NUM_WRITE-1:0] WDATA
);
   reg [DW-1:0] regfile [(1<<AW)-1:0];
   reg [DW-1:0] ff_dout [NUM_READ-1:0];
   genvar i;
   integer j;
   always @(posedge CLK)
      for(j=0;j<NUM_WRITE;j=j+1) 
         if (WE[j])
            regfile[WADDR[j*AW +: AW]] <= WDATA[j*DW +: DW];
   generate
      for(i=0;i<NUM_READ;i=i+1)
         begin
            always @(posedge CLK)
               if (RE[i])
                  ff_dout[i] <= regfile[RADDR[i*AW +: AW]];
            assign RDATA[i*DW +: DW] = ff_dout[i];
         end
   endgenerate
endmodule
module ysyx_20210479
(
   input	clock,
   input	reset,
   input	io_interrupt,
   input io_master_awready,
   output io_master_awvalid,
   output [31:0]	io_master_awaddr,
   output [3:0]	io_master_awid,
   output [7:0]	io_master_awlen,
   output [2:0]	io_master_awsize,
   output [1:0]	io_master_awburst,
   input io_master_wready,
   output io_master_wvalid,
   output [63:0]	io_master_wdata,
   output [7:0]	io_master_wstrb,
   output io_master_wlast,
   output io_master_bready,
   input io_master_bvalid,
   input	[1:0]	io_master_bresp,
   input	[3:0]	io_master_bid,
   input io_master_arready,
   output io_master_arvalid,
   output [31:0]	io_master_araddr,
   output [3:0]	io_master_arid,
   output [7:0]	io_master_arlen,
   output [2:0]	io_master_arsize,
   output io_master_rready,
   input io_master_rvalid,
   input	[1:0]	io_master_rresp,
   input	[63:0]	io_master_rdata,
   input io_master_rlast,
   input	[3:0]	io_master_rid,
   output io_slave_awready,
	input io_slave_awvalid,
	input	[31:0]	io_slave_awaddr,
	input	[3:0]	io_slave_awid,
	input	[7:0]	io_slave_awlen,
	input	[2:0]	io_slave_awsize,
	input	[1:0]	io_slave_awburst,
	output io_slave_wready,
   input io_slave_wvalid,
	input	[63:0]	io_slave_wdata,
	input	[7:0]	io_slave_wstrb,
	input io_slave_wlast,
	input io_slave_bready,
	output io_slave_bvalid,
	output [1:0]	io_slave_bresp,
	output [3:0]	io_slave_bid,
	output io_slave_arready,
	input io_slave_arvalid,
	input	[31:0]	io_slave_araddr,
	input	[3:0]	io_slave_arid,
	input	[7:0]	io_slave_arlen,
	input	[2:0]	io_slave_arsize,
   output [1:0]	io_master_arburst,
	input	[1:0]	io_slave_arburst,
	input io_slave_rready,
	output io_slave_rvalid,
	output [1:0]	io_slave_rresp,
	output [63:0]	io_slave_rdata,
	output io_slave_rlast,
	output [3:0]	io_slave_rid
);
   localparam                           CONFIG_AW = 32;
   localparam                           CONFIG_DW = 32;
   localparam                           CONFIG_P_DW = 5;
   localparam                           CONFIG_P_FETCH_WIDTH = 1;
   localparam                           CONFIG_P_ISSUE_WIDTH = 1;
   localparam                           CONFIG_P_PAGE_SIZE = 13;
   localparam                           CONFIG_IC_P_LINE = 6;
   localparam                           CONFIG_IC_P_SETS = 4;
   localparam                           CONFIG_IC_P_WAYS = 1;
   localparam                           CONFIG_DC_P_LINE = 6;
   localparam                           CONFIG_DC_P_SETS = 4;
   localparam                           CONFIG_DC_P_WAYS = 1;
   localparam                           CONFIG_PHT_P_NUM = 2;
   localparam                           CONFIG_BTB_P_NUM = 2;
   localparam                           CONFIG_P_IQ_DEPTH = 2;
   localparam                           CONFIG_ENABLE_MUL = 0;
   localparam                           CONFIG_ENABLE_DIV = 0;
   localparam                           CONFIG_ENABLE_DIVU = 0;
   localparam                           CONFIG_ENABLE_MOD = 0;
   localparam                           CONFIG_ENABLE_MODU = 0;
   localparam                           CONFIG_ENABLE_ASR = 1;
   localparam                           CONFIG_IMMU_ENABLE_UNCACHED_SEG = 1;
   localparam                           CONFIG_DMMU_ENABLE_UNCACHED_SEG = 1;
   localparam                           CONFIG_DTLB_P_SETS = 7;
   localparam                           CONFIG_ITLB_P_SETS = 7;
   localparam [CONFIG_AW-1:0]           CONFIG_ERST_VECTOR = 32'h80000000; 
   localparam [CONFIG_AW-1:0]           CONFIG_EITM_VECTOR = 32'h80000000 + 32'h1c;
   localparam [CONFIG_AW-1:0]           CONFIG_EIPF_VECTOR = 32'h80000000 + 32'h14;
   localparam [CONFIG_AW-1:0]           CONFIG_ESYSCALL_VECTOR = 32'h80000000 + 32'hc;
   localparam [CONFIG_AW-1:0]           CONFIG_EINSN_VECTOR = 32'h80000000 + 32'h4;
   localparam [CONFIG_AW-1:0]           CONFIG_EIRQ_VECTOR = 32'h80000000 + 32'h8;
   localparam [CONFIG_AW-1:0]           CONFIG_EDTM_VECTOR = 32'h80000000 + 32'h20;
   localparam [CONFIG_AW-1:0]           CONFIG_EDPF_VECTOR = 32'h80000000 + 32'h18;
   localparam [CONFIG_AW-1:0]           CONFIG_EALIGN_VECTOR = 32'h80000000 + 32'h24;
   localparam                           CONFIG_NUM_IRQ = 32;
   localparam AXI_P_DW_BYTES   = 3; 
   localparam AXI_UNCACHED_P_DW_BYTES = 2; 
   localparam AXI_ADDR_WIDTH    = 32;
   localparam AXI_ID_WIDTH      = 4;
   localparam AXI_USER_WIDTH    = 1;
   wire [AXI_ADDR_WIDTH-1:0] dbus_ARADDR;       
   wire [1:0]           dbus_ARBURST;           
   wire [3:0]           dbus_ARCACHE;           
   wire [AXI_ID_WIDTH-1:0] dbus_ARID;           
   wire [7:0]           dbus_ARLEN;             
   wire                 dbus_ARLOCK;            
   wire [2:0]           dbus_ARPROT;            
   wire [3:0]           dbus_ARQOS;             
   wire                 dbus_ARREADY;           
   wire [3:0]           dbus_ARREGION;          
   wire [2:0]           dbus_ARSIZE;            
   wire [AXI_USER_WIDTH-1:0] dbus_ARUSER;       
   wire                 dbus_ARVALID;           
   wire [AXI_ADDR_WIDTH-1:0] dbus_AWADDR;       
   wire [1:0]           dbus_AWBURST;           
   wire [3:0]           dbus_AWCACHE;           
   wire [AXI_ID_WIDTH-1:0] dbus_AWID;           
   wire [7:0]           dbus_AWLEN;             
   wire                 dbus_AWLOCK;            
   wire [2:0]           dbus_AWPROT;            
   wire [3:0]           dbus_AWQOS;             
   wire                 dbus_AWREADY;           
   wire [3:0]           dbus_AWREGION;          
   wire [2:0]           dbus_AWSIZE;            
   wire [AXI_USER_WIDTH-1:0] dbus_AWUSER;       
   wire                 dbus_AWVALID;           
   wire [AXI_ID_WIDTH-1:0] dbus_BID;            
   wire                 dbus_BREADY;            
   wire [1:0]           dbus_BRESP;             
   wire [AXI_USER_WIDTH-1:0] dbus_BUSER;        
   wire                 dbus_BVALID;            
   wire [(1<<AXI_P_DW_BYTES)*8-1:0] dbus_RDATA; 
   wire [AXI_ID_WIDTH-1:0] dbus_RID;            
   wire                 dbus_RLAST;             
   wire                 dbus_RREADY;            
   wire [1:0]           dbus_RRESP;             
   wire [AXI_USER_WIDTH-1:0] dbus_RUSER;        
   wire                 dbus_RVALID;            
   wire [(1<<AXI_P_DW_BYTES)*8-1:0] dbus_WDATA; 
   wire                 dbus_WLAST;             
   wire                 dbus_WREADY;            
   wire [(1<<AXI_P_DW_BYTES)-1:0] dbus_WSTRB;   
   wire [AXI_USER_WIDTH-1:0] dbus_WUSER;        
   wire                 dbus_WVALID;            
   wire [AXI_ADDR_WIDTH-1:0] ibus_ARADDR;       
   wire [1:0]           ibus_ARBURST;           
   wire [3:0]           ibus_ARCACHE;           
   wire [AXI_ID_WIDTH-1:0] ibus_ARID;           
   wire [7:0]           ibus_ARLEN;             
   wire                 ibus_ARLOCK;            
   wire [2:0]           ibus_ARPROT;            
   wire [3:0]           ibus_ARQOS;             
   wire                 ibus_ARREADY;           
   wire [3:0]           ibus_ARREGION;          
   wire [2:0]           ibus_ARSIZE;            
   wire [AXI_USER_WIDTH-1:0] ibus_ARUSER;       
   wire                 ibus_ARVALID;           
   wire                 ibus_AWREADY;           
   wire [AXI_ID_WIDTH-1:0] ibus_BID;            
   wire [1:0]           ibus_BRESP;             
   wire [AXI_USER_WIDTH-1:0] ibus_BUSER;        
   wire                 ibus_BVALID;            
   wire [(1<<AXI_P_DW_BYTES)*8-1:0] ibus_RDATA; 
   wire [AXI_ID_WIDTH-1:0] ibus_RID;            
   wire                 ibus_RLAST;             
   wire                 ibus_RREADY;            
   wire [1:0]           ibus_RRESP;             
   wire [AXI_USER_WIDTH-1:0] ibus_RUSER;        
   wire                 ibus_RVALID;            
   wire                 ibus_WREADY;            
   wire                 tsc_irq;                
   wire [3:0]           io_master_arcache;      
   wire                 io_master_arlock;       
   wire [2:0]           io_master_arprot;       
   wire [3:0]           io_master_arqos;        
   wire [3:0]           io_master_arregion;     
   wire [AXI_USER_WIDTH-1:0] io_master_aruser;  
   wire [3:0]           io_master_awcache;      
   wire                 io_master_awlock;       
   wire [2:0]           io_master_awprot;       
   wire [3:0]           io_master_awqos;        
   wire [3:0]           io_master_awregion;     
   wire [AXI_USER_WIDTH-1:0] io_master_awuser;  
   wire [AXI_USER_WIDTH-1:0] io_master_wuser;   
   wire                 clk;                    
   wire                 rst;                    
   wire  [CONFIG_NUM_IRQ-1:0] irqs;             
   wire  [AXI_ADDR_WIDTH-1:0] ibus_AWADDR;      
   wire  [1:0]          ibus_AWBURST;           
   wire  [3:0]          ibus_AWCACHE;           
   wire  [AXI_ID_WIDTH-1:0] ibus_AWID;          
   wire  [7:0]          ibus_AWLEN;             
   wire                 ibus_AWLOCK;            
   wire  [2:0]          ibus_AWPROT;            
   wire  [3:0]          ibus_AWQOS;             
   wire  [3:0]          ibus_AWREGION;          
   wire  [2:0]          ibus_AWSIZE;            
   wire  [AXI_USER_WIDTH-1:0] ibus_AWUSER;      
   wire                 ibus_AWVALID;           
   wire                 ibus_BREADY;            
   wire  [(1<<AXI_P_DW_BYTES)*8-1:0] ibus_WDATA;
   wire                 ibus_WLAST;             
   wire  [(1<<AXI_P_DW_BYTES)-1:0] ibus_WSTRB;  
   wire  [AXI_USER_WIDTH-1:0] ibus_WUSER;       
   wire                 ibus_WVALID;            
   wire  [AXI_USER_WIDTH-1:0] io_master_buser;  
   wire  [AXI_USER_WIDTH-1:0] io_master_ruser;  
   assign clk = clock;
   assign rst = reset;
   ysyx_20210479_ncpu64k
      #(
        .CONFIG_AW                      (CONFIG_AW),
        .CONFIG_DW                      (CONFIG_DW),
        .CONFIG_P_DW                    (CONFIG_P_DW),
        .CONFIG_P_FETCH_WIDTH           (CONFIG_P_FETCH_WIDTH),
        .CONFIG_P_ISSUE_WIDTH           (CONFIG_P_ISSUE_WIDTH),
        .CONFIG_P_PAGE_SIZE             (CONFIG_P_PAGE_SIZE),
        .CONFIG_IC_P_LINE               (CONFIG_IC_P_LINE),
        .CONFIG_IC_P_SETS               (CONFIG_IC_P_SETS),
        .CONFIG_IC_P_WAYS               (CONFIG_IC_P_WAYS),
        .CONFIG_DC_P_LINE               (CONFIG_DC_P_LINE),
        .CONFIG_DC_P_SETS               (CONFIG_DC_P_SETS),
        .CONFIG_DC_P_WAYS               (CONFIG_DC_P_WAYS),
        .CONFIG_PHT_P_NUM               (CONFIG_PHT_P_NUM),
        .CONFIG_BTB_P_NUM               (CONFIG_BTB_P_NUM),
        .CONFIG_P_IQ_DEPTH              (CONFIG_P_IQ_DEPTH),
        .CONFIG_ENABLE_MUL              (CONFIG_ENABLE_MUL),
        .CONFIG_ENABLE_DIV              (CONFIG_ENABLE_DIV),
        .CONFIG_ENABLE_DIVU             (CONFIG_ENABLE_DIVU),
        .CONFIG_ENABLE_MOD              (CONFIG_ENABLE_MOD),
        .CONFIG_ENABLE_MODU             (CONFIG_ENABLE_MODU),
        .CONFIG_ENABLE_ASR              (CONFIG_ENABLE_ASR),
        .CONFIG_IMMU_ENABLE_UNCACHED_SEG(CONFIG_IMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_DMMU_ENABLE_UNCACHED_SEG(CONFIG_DMMU_ENABLE_UNCACHED_SEG),
        .CONFIG_DTLB_P_SETS             (CONFIG_DTLB_P_SETS),
        .CONFIG_ITLB_P_SETS             (CONFIG_ITLB_P_SETS),
        .CONFIG_ERST_VECTOR             (CONFIG_ERST_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EITM_VECTOR             (CONFIG_EITM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIPF_VECTOR             (CONFIG_EIPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_ESYSCALL_VECTOR         (CONFIG_ESYSCALL_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EINSN_VECTOR            (CONFIG_EINSN_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EIRQ_VECTOR             (CONFIG_EIRQ_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDTM_VECTOR             (CONFIG_EDTM_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EDPF_VECTOR             (CONFIG_EDPF_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_EALIGN_VECTOR           (CONFIG_EALIGN_VECTOR[CONFIG_AW-1:0]),
        .CONFIG_NUM_IRQ                 (CONFIG_NUM_IRQ),
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_UNCACHED_P_DW_BYTES        (AXI_UNCACHED_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_CORE
      (
       .ibus_ARVALID                    (ibus_ARVALID),
       .ibus_ARADDR                     (ibus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .ibus_ARPROT                     (ibus_ARPROT[2:0]),
       .ibus_ARID                       (ibus_ARID[AXI_ID_WIDTH-1:0]),
       .ibus_ARUSER                     (ibus_ARUSER[AXI_USER_WIDTH-1:0]),
       .ibus_ARLEN                      (ibus_ARLEN[7:0]),
       .ibus_ARSIZE                     (ibus_ARSIZE[2:0]),
       .ibus_ARBURST                    (ibus_ARBURST[1:0]),
       .ibus_ARLOCK                     (ibus_ARLOCK),
       .ibus_ARCACHE                    (ibus_ARCACHE[3:0]),
       .ibus_ARQOS                      (ibus_ARQOS[3:0]),
       .ibus_ARREGION                   (ibus_ARREGION[3:0]),
       .ibus_RREADY                     (ibus_RREADY),
       .dbus_ARVALID                    (dbus_ARVALID),
       .dbus_ARADDR                     (dbus_ARADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_ARPROT                     (dbus_ARPROT[2:0]),
       .dbus_ARID                       (dbus_ARID[AXI_ID_WIDTH-1:0]),
       .dbus_ARUSER                     (dbus_ARUSER[AXI_USER_WIDTH-1:0]),
       .dbus_ARLEN                      (dbus_ARLEN[7:0]),
       .dbus_ARSIZE                     (dbus_ARSIZE[2:0]),
       .dbus_ARBURST                    (dbus_ARBURST[1:0]),
       .dbus_ARLOCK                     (dbus_ARLOCK),
       .dbus_ARCACHE                    (dbus_ARCACHE[3:0]),
       .dbus_ARQOS                      (dbus_ARQOS[3:0]),
       .dbus_ARREGION                   (dbus_ARREGION[3:0]),
       .dbus_RREADY                     (dbus_RREADY),
       .dbus_AWVALID                    (dbus_AWVALID),
       .dbus_AWADDR                     (dbus_AWADDR[AXI_ADDR_WIDTH-1:0]),
       .dbus_AWPROT                     (dbus_AWPROT[2:0]),
       .dbus_AWID                       (dbus_AWID[AXI_ID_WIDTH-1:0]),
       .dbus_AWUSER                     (dbus_AWUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWLEN                      (dbus_AWLEN[7:0]),
       .dbus_AWSIZE                     (dbus_AWSIZE[2:0]),
       .dbus_AWBURST                    (dbus_AWBURST[1:0]),
       .dbus_AWLOCK                     (dbus_AWLOCK),
       .dbus_AWCACHE                    (dbus_AWCACHE[3:0]),
       .dbus_AWQOS                      (dbus_AWQOS[3:0]),
       .dbus_AWREGION                   (dbus_AWREGION[3:0]),
       .dbus_WVALID                     (dbus_WVALID),
       .dbus_WDATA                      (dbus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_WSTRB                      (dbus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]),
       .dbus_WLAST                      (dbus_WLAST),
       .dbus_WUSER                      (dbus_WUSER[AXI_USER_WIDTH-1:0]),
       .dbus_BREADY                     (dbus_BREADY),
       .tsc_irq                         (tsc_irq),
       .clk                             (clk),
       .rst                             (rst),
       .ibus_ARREADY                    (ibus_ARREADY),
       .ibus_RVALID                     (ibus_RVALID),
       .ibus_RDATA                      (ibus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .ibus_RLAST                      (ibus_RLAST),
       .ibus_RRESP                      (ibus_RRESP[1:0]),
       .ibus_RID                        (ibus_RID[AXI_ID_WIDTH-1:0]),
       .ibus_RUSER                      (ibus_RUSER[AXI_USER_WIDTH-1:0]),
       .dbus_ARREADY                    (dbus_ARREADY),
       .dbus_RVALID                     (dbus_RVALID),
       .dbus_RDATA                      (dbus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]),
       .dbus_RRESP                      (dbus_RRESP[1:0]),
       .dbus_RLAST                      (dbus_RLAST),
       .dbus_RID                        (dbus_RID[AXI_ID_WIDTH-1:0]),
       .dbus_RUSER                      (dbus_RUSER[AXI_USER_WIDTH-1:0]),
       .dbus_AWREADY                    (dbus_AWREADY),
       .dbus_WREADY                     (dbus_WREADY),
       .dbus_BVALID                     (dbus_BVALID),
       .dbus_BRESP                      (dbus_BRESP[1:0]),
       .dbus_BID                        (dbus_BID[AXI_ID_WIDTH-1:0]),
       .dbus_BUSER                      (dbus_BUSER[AXI_USER_WIDTH-1:0]),
       .irqs                            (irqs[CONFIG_NUM_IRQ-1:0]));
   axi4_arbiter
      #(
        .AXI_P_DW_BYTES                 (AXI_P_DW_BYTES),
        .AXI_ADDR_WIDTH                 (AXI_ADDR_WIDTH),
        .AXI_ID_WIDTH                   (AXI_ID_WIDTH),
        .AXI_USER_WIDTH                 (AXI_USER_WIDTH))
   U_AXI4_ARBITER
      (
       .s0_ARREADY                      (ibus_ARREADY),          
       .s0_RVALID                       (ibus_RVALID),           
       .s0_RDATA                        (ibus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .s0_RRESP                        (ibus_RRESP[1:0]),       
       .s0_RLAST                        (ibus_RLAST),            
       .s0_RID                          (ibus_RID[AXI_ID_WIDTH-1:0]), 
       .s0_RUSER                        (ibus_RUSER[AXI_USER_WIDTH-1:0]), 
       .s0_AWREADY                      (ibus_AWREADY),          
       .s0_WREADY                       (ibus_WREADY),           
       .s0_BVALID                       (ibus_BVALID),           
       .s0_BRESP                        (ibus_BRESP[1:0]),       
       .s0_BID                          (ibus_BID[AXI_ID_WIDTH-1:0]), 
       .s0_BUSER                        (ibus_BUSER[AXI_USER_WIDTH-1:0]), 
       .s1_ARREADY                      (dbus_ARREADY),          
       .s1_RVALID                       (dbus_RVALID),           
       .s1_RDATA                        (dbus_RDATA[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .s1_RRESP                        (dbus_RRESP[1:0]),       
       .s1_RLAST                        (dbus_RLAST),            
       .s1_RID                          (dbus_RID[AXI_ID_WIDTH-1:0]), 
       .s1_RUSER                        (dbus_RUSER[AXI_USER_WIDTH-1:0]), 
       .s1_AWREADY                      (dbus_AWREADY),          
       .s1_WREADY                       (dbus_WREADY),           
       .s1_BVALID                       (dbus_BVALID),           
       .s1_BRESP                        (dbus_BRESP[1:0]),       
       .s1_BID                          (dbus_BID[AXI_ID_WIDTH-1:0]), 
       .s1_BUSER                        (dbus_BUSER[AXI_USER_WIDTH-1:0]), 
       .m_ARVALID                       (io_master_arvalid),     
       .m_ARADDR                        (io_master_araddr[AXI_ADDR_WIDTH-1:0]), 
       .m_ARPROT                        (io_master_arprot[2:0]), 
       .m_ARID                          (io_master_arid[AXI_ID_WIDTH-1:0]), 
       .m_ARUSER                        (io_master_aruser[AXI_USER_WIDTH-1:0]), 
       .m_ARLEN                         (io_master_arlen[7:0]),  
       .m_ARSIZE                        (io_master_arsize[2:0]), 
       .m_ARBURST                       (io_master_arburst[1:0]), 
       .m_ARLOCK                        (io_master_arlock),      
       .m_ARCACHE                       (io_master_arcache[3:0]), 
       .m_ARQOS                         (io_master_arqos[3:0]),  
       .m_ARREGION                      (io_master_arregion[3:0]), 
       .m_RREADY                        (io_master_rready),      
       .m_AWVALID                       (io_master_awvalid),     
       .m_AWADDR                        (io_master_awaddr[AXI_ADDR_WIDTH-1:0]), 
       .m_AWPROT                        (io_master_awprot[2:0]), 
       .m_AWID                          (io_master_awid[AXI_ID_WIDTH-1:0]), 
       .m_AWUSER                        (io_master_awuser[AXI_USER_WIDTH-1:0]), 
       .m_AWLEN                         (io_master_awlen[7:0]),  
       .m_AWSIZE                        (io_master_awsize[2:0]), 
       .m_AWBURST                       (io_master_awburst[1:0]), 
       .m_AWLOCK                        (io_master_awlock),      
       .m_AWCACHE                       (io_master_awcache[3:0]), 
       .m_AWQOS                         (io_master_awqos[3:0]),  
       .m_AWREGION                      (io_master_awregion[3:0]), 
       .m_WVALID                        (io_master_wvalid),      
       .m_WDATA                         (io_master_wdata[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .m_WSTRB                         (io_master_wstrb[(1<<AXI_P_DW_BYTES)-1:0]), 
       .m_WLAST                         (io_master_wlast),       
       .m_WUSER                         (io_master_wuser[AXI_USER_WIDTH-1:0]), 
       .m_BREADY                        (io_master_bready),      
       .clk                             (clk),
       .rst                             (rst),
       .s0_ARVALID                      (ibus_ARVALID),          
       .s0_ARADDR                       (ibus_ARADDR[AXI_ADDR_WIDTH-1:0]), 
       .s0_ARPROT                       (ibus_ARPROT[2:0]),      
       .s0_ARID                         (ibus_ARID[AXI_ID_WIDTH-1:0]), 
       .s0_ARUSER                       (ibus_ARUSER[AXI_USER_WIDTH-1:0]), 
       .s0_ARLEN                        (ibus_ARLEN[7:0]),       
       .s0_ARSIZE                       (ibus_ARSIZE[2:0]),      
       .s0_ARBURST                      (ibus_ARBURST[1:0]),     
       .s0_ARLOCK                       (ibus_ARLOCK),           
       .s0_ARCACHE                      (ibus_ARCACHE[3:0]),     
       .s0_ARQOS                        (ibus_ARQOS[3:0]),       
       .s0_ARREGION                     (ibus_ARREGION[3:0]),    
       .s0_RREADY                       (ibus_RREADY),           
       .s0_AWVALID                      (ibus_AWVALID),          
       .s0_AWADDR                       (ibus_AWADDR[AXI_ADDR_WIDTH-1:0]), 
       .s0_AWPROT                       (ibus_AWPROT[2:0]),      
       .s0_AWID                         (ibus_AWID[AXI_ID_WIDTH-1:0]), 
       .s0_AWUSER                       (ibus_AWUSER[AXI_USER_WIDTH-1:0]), 
       .s0_AWLEN                        (ibus_AWLEN[7:0]),       
       .s0_AWSIZE                       (ibus_AWSIZE[2:0]),      
       .s0_AWBURST                      (ibus_AWBURST[1:0]),     
       .s0_AWLOCK                       (ibus_AWLOCK),           
       .s0_AWCACHE                      (ibus_AWCACHE[3:0]),     
       .s0_AWQOS                        (ibus_AWQOS[3:0]),       
       .s0_AWREGION                     (ibus_AWREGION[3:0]),    
       .s0_WVALID                       (ibus_WVALID),           
       .s0_WDATA                        (ibus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .s0_WSTRB                        (ibus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]), 
       .s0_WLAST                        (ibus_WLAST),            
       .s0_WUSER                        (ibus_WUSER[AXI_USER_WIDTH-1:0]), 
       .s0_BREADY                       (ibus_BREADY),           
       .s1_ARVALID                      (dbus_ARVALID),          
       .s1_ARADDR                       (dbus_ARADDR[AXI_ADDR_WIDTH-1:0]), 
       .s1_ARPROT                       (dbus_ARPROT[2:0]),      
       .s1_ARID                         (dbus_ARID[AXI_ID_WIDTH-1:0]), 
       .s1_ARUSER                       (dbus_ARUSER[AXI_USER_WIDTH-1:0]), 
       .s1_ARLEN                        (dbus_ARLEN[7:0]),       
       .s1_ARSIZE                       (dbus_ARSIZE[2:0]),      
       .s1_ARBURST                      (dbus_ARBURST[1:0]),     
       .s1_ARLOCK                       (dbus_ARLOCK),           
       .s1_ARCACHE                      (dbus_ARCACHE[3:0]),     
       .s1_ARQOS                        (dbus_ARQOS[3:0]),       
       .s1_ARREGION                     (dbus_ARREGION[3:0]),    
       .s1_RREADY                       (dbus_RREADY),           
       .s1_AWVALID                      (dbus_AWVALID),          
       .s1_AWADDR                       (dbus_AWADDR[AXI_ADDR_WIDTH-1:0]), 
       .s1_AWPROT                       (dbus_AWPROT[2:0]),      
       .s1_AWID                         (dbus_AWID[AXI_ID_WIDTH-1:0]), 
       .s1_AWUSER                       (dbus_AWUSER[AXI_USER_WIDTH-1:0]), 
       .s1_AWLEN                        (dbus_AWLEN[7:0]),       
       .s1_AWSIZE                       (dbus_AWSIZE[2:0]),      
       .s1_AWBURST                      (dbus_AWBURST[1:0]),     
       .s1_AWLOCK                       (dbus_AWLOCK),           
       .s1_AWCACHE                      (dbus_AWCACHE[3:0]),     
       .s1_AWQOS                        (dbus_AWQOS[3:0]),       
       .s1_AWREGION                     (dbus_AWREGION[3:0]),    
       .s1_WVALID                       (dbus_WVALID),           
       .s1_WDATA                        (dbus_WDATA[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .s1_WSTRB                        (dbus_WSTRB[(1<<AXI_P_DW_BYTES)-1:0]), 
       .s1_WLAST                        (dbus_WLAST),            
       .s1_WUSER                        (dbus_WUSER[AXI_USER_WIDTH-1:0]), 
       .s1_BREADY                       (dbus_BREADY),           
       .m_ARREADY                       (io_master_arready),     
       .m_RVALID                        (io_master_rvalid),      
       .m_RDATA                         (io_master_rdata[(1<<AXI_P_DW_BYTES)*8-1:0]), 
       .m_RRESP                         (io_master_rresp[1:0]),  
       .m_RLAST                         (io_master_rlast),       
       .m_RID                           (io_master_rid[AXI_ID_WIDTH-1:0]), 
       .m_RUSER                         (io_master_ruser[AXI_USER_WIDTH-1:0]), 
       .m_AWREADY                       (io_master_awready),     
       .m_WREADY                        (io_master_wready),      
       .m_BVALID                        (io_master_bvalid),      
       .m_BRESP                         (io_master_bresp[1:0]),  
       .m_BID                           (io_master_bid[AXI_ID_WIDTH-1:0]), 
       .m_BUSER                         (io_master_buser[AXI_USER_WIDTH-1:0])); 
   assign ibus_AWADDR = 'b0;
   assign ibus_AWBURST = 'b0;
   assign ibus_AWCACHE = 'b0;
   assign ibus_AWID = 'b0;
   assign ibus_AWLEN = 'b0;
   assign ibus_AWLOCK = 'b0;
   assign ibus_AWPROT = 'b0;
   assign ibus_AWQOS = 'b0;
   assign ibus_AWREGION = 'b0;
   assign ibus_AWSIZE = 'b0;
   assign ibus_AWUSER = 'b0;
   assign ibus_AWVALID = 'b0;
   assign ibus_BREADY = 'b0;
   assign ibus_WDATA = 'b0;
   assign ibus_WLAST = 'b0;
   assign ibus_WSTRB = 'b0;
   assign ibus_WUSER = 'b0;
   assign ibus_WVALID = 'b0;
   assign io_master_buser = 'b0;
   assign io_master_ruser = 'b0;
   assign irqs[0] = tsc_irq;
   assign irqs[30:1] = 'b0;
   assign irqs[31] = io_interrupt;
   assign io_slave_awready = 'b0;
	assign io_slave_wready = 'b0;
	assign io_slave_bvalid = 'b0;
	assign io_slave_bresp = 'b0;
	assign io_slave_bid = 'b0;
	assign io_slave_arready = 'b0;
	assign io_slave_rvalid = 'b0;
	assign io_slave_rresp = 'b0;
	assign io_slave_rdata = 'b0;
	assign io_slave_rlast = 'b0;
	assign io_slave_rid = 'b0;
endmodule
